`timescale 1ns/1ps

module ND6( o, i0, i1, i2, i3, i4, i5 );
    input  i0, i1, i2, i3, i4, i5;
    output o;
    wire   dummy0, dummy1;
    ND3 nd0( dummy0, i0, i1, i2 );
    ND3 nd1( dummy1, i3, i4, i5 );
    OR2 ret( o, dummy0, dummy1 );
endmodule

module OR6( o, i0, i1, i2, i3, i4, i5 );
    input  i0, i1, i2, i3, i4, i5;
    output o;
    wire   dummy;
    OR4 or_( dummy, i0, i1, i2, i3 );
    OR3 ret( o, i4, i5, dummy );
endmodule

module AN6( o, i0, i1, i2, i3, i4, i5 );
    input  i0, i1, i2, i3, i4, i5;
    output o;
    wire   dummy;
    AN4 an_( dummy, i0, i1, i2, i3 );
    AN3 ret( o, i4, i5, dummy );
endmodule

module OR5( o, i0, i1, i2, i3, i4 );
    input  i0, i1, i2, i3, i4;
    output o;
    wire   dummy;
    OR3 or_( dummy, i0, i1, i2 );
    OR3 ret( o, i3, i4, dummy );
endmodule

module AN5( o, i0, i1, i2, i3, i4 );
    input  i0, i1, i2, i3, i4;
    output o;
    wire   dummy;
    AN3 an_( dummy, i0, i1, i2 );
    AN3 ret( o, i3, i4, dummy );
endmodule

module foobar( o, A, B );
    input  A, B;
    output o;
    wire   a;
    IV  inv( a, A );
    AN2 ret( o, a, B );
endmodule

module OR15( o, i );
    input [14:0] i;
    output       o;
    wire dummy0, dummy1, dummy2, dummy3;
    OR4 or_0_3( dummy0, i[0],   i[1],   i[2],   i[3]   );
    OR4 or_4_7( dummy1, i[4],   i[5],   i[6],   i[7]   );
    OR4 or_8_B( dummy2, i[8],   i[9],   i[10],  i[11]  );
    OR3 or_C_E( dummy3, i[12],  i[13],  i[14]          );
    OR4 ret   ( o,      dummy0, dummy1, dummy2, dummy3 );
endmodule

module OR20( o, i );
    input  [19:0] i;
    output        o;
    wire   [5:0]  dummy;
    OR4 or_0_3( dummy[0], i[0],     i[1],     i[2],     i[3]   );
    OR4 or_4_7( dummy[1], i[4],     i[5],     i[6],     i[7]   );
    OR4 or_8_B( dummy[2], i[8],     i[9],     i[10],    i[11]  );
    OR4 or_C_F( dummy[3], i[12],    i[13],    i[14],    i[15]  );
    OR4 or_G_J( dummy[4], i[16],    i[17],    i[18],    i[19]  );
    OR4 or_0_F( dummy[5], dummy[0], dummy[1], dummy[2], dummy[3] );
    OR2 ret   ( o       , dummy[5], dummy[4] );
endmodule

module OR32( o, i );
    input  [31:0] i;
    output        o;
    wire   [9:0]  dummy;
    OR4 or_0_3( dummy[0], i[0],     i[1],     i[2],     i[3]   );
    OR4 or_4_7( dummy[1], i[4],     i[5],     i[6],     i[7]   );
    OR4 or_8_B( dummy[2], i[8],     i[9],     i[10],    i[11]  );
    OR4 or_C_F( dummy[3], i[12],    i[13],    i[14],    i[15]  );
    OR4 or_G_J( dummy[4], i[16],    i[17],    i[18],    i[19]  );
    OR4 or_K_N( dummy[5], i[20],    i[21],    i[22],    i[23]  );
    OR4 or_O_R( dummy[6], i[24],    i[25],    i[26],    i[27]  );
    OR4 or_S_V( dummy[7], i[28],    i[29],    i[30],    i[31]  );
    OR4 or_0_F( dummy[8], dummy[0], dummy[1], dummy[2], dummy[3] );
    OR4 or_G_V( dummy[9], dummy[4], dummy[5], dummy[6], dummy[7] );
    OR2 ret   ( o       , dummy[8], dummy[9] );
endmodule

module AN64( o, i );
    input  [63:0] i;
    output        o;
    wire   [19:0]  dummy;
    AN4 or_00  ( dummy[ 0], i[0],      i[1],      i[2],      i[3]      );
    AN4 or_01  ( dummy[ 1], i[4],      i[5],      i[6],      i[7]      );
    AN4 or_02  ( dummy[ 2], i[8],      i[9],      i[10],     i[11]     );
    AN4 or_03  ( dummy[ 3], i[12],     i[13],     i[14],     i[15]     );
    AN4 or_04  ( dummy[ 4], i[16],     i[17],     i[18],     i[19]     );
    AN4 or_05  ( dummy[ 5], i[20],     i[21],     i[22],     i[23]     );
    AN4 or_06  ( dummy[ 6], i[24],     i[25],     i[26],     i[27]     );
    AN4 or_07  ( dummy[ 7], i[28],     i[29],     i[30],     i[31]     );
    AN4 or_08  ( dummy[ 8], i[32],     i[33],     i[34],     i[35]     );
    AN4 or_09  ( dummy[ 9], i[36],     i[37],     i[38],     i[39]     );
    AN4 or_10  ( dummy[10], i[40],     i[41],     i[42],     i[43]     );
    AN4 or_11  ( dummy[11], i[44],     i[45],     i[46],     i[47]     );
    AN4 or_12  ( dummy[12], i[48],     i[49],     i[50],     i[51]     );
    AN4 or_13  ( dummy[13], i[52],     i[53],     i[54],     i[55]     );
    AN4 or_14  ( dummy[14], i[56],     i[57],     i[58],     i[59]     );
    AN4 or_15  ( dummy[15], i[60],     i[61],     i[62],     i[63]     );
    AN4 d_00_03( dummy[16], dummy[0],  dummy[1],  dummy[2],  dummy[3]  );
    AN4 d_04_07( dummy[17], dummy[4],  dummy[5],  dummy[6],  dummy[7]  );
    AN4 d_08_11( dummy[18], dummy[8],  dummy[9],  dummy[10], dummy[11] );
    AN4 d_12_15( dummy[19], dummy[12], dummy[13], dummy[14], dummy[15] );
    AN4 ret    ( o,         dummy[16], dummy[17], dummy[18], dummy[19] );
endmodule

`define wires_2_6 \
    wire  AB, AC, AD, AE, AF, BC, BD, BE, BF, CD, CE, CF, DE, DF, EF; \
    AN2 gate_AB ( AB, A, B ); \
    AN2 gate_AC ( AC, A, C ); \
    AN2 gate_AD ( AD, A, D ); \
    AN2 gate_AE ( AE, A, E ); \
    AN2 gate_AF ( AF, A, F ); \
    AN2 gate_BC ( BC, B, C ); \
    AN2 gate_BD ( BD, B, D ); \
    AN2 gate_BE ( BE, B, E ); \
    AN2 gate_BF ( BF, B, F ); \
    AN2 gate_CD ( CD, C, D ); \
    AN2 gate_CE ( CE, C, E ); \
    AN2 gate_CF ( CF, C, F ); \
    AN2 gate_DE ( DE, D, E ); \
    AN2 gate_DF ( DF, D, F ); \
    AN2 gate_EF ( EF, E, F );

`define wires_3_6 \
    wire  ABC, ABD, ABE, ABF, ACD, ACE, ACF, ADE, ADF, AEF, BCD, BCE, BCF, BDE, BDF, BEF, CDE, CDF, CEF, DEF; \
    AN3 gate_ABC( ABC, A, B, C ); \
    AN3 gate_ABD( ABD, A, B, D ); \
    AN3 gate_ABE( ABE, A, B, E ); \
    AN3 gate_ABF( ABF, A, B, F ); \
    AN3 gate_ACD( ACD, A, C, D ); \
    AN3 gate_ACE( ACE, A, C, E ); \
    AN3 gate_ACF( ACF, A, C, F ); \
    AN3 gate_ADE( ADE, A, D, E ); \
    AN3 gate_ADF( ADF, A, D, F ); \
    AN3 gate_AEF( AEF, A, E, F ); \
    AN3 gate_BCD( BCD, B, C, D ); \
    AN3 gate_BCE( BCE, B, C, E ); \
    AN3 gate_BCF( BCF, B, C, F ); \
    AN3 gate_BDE( BDE, B, D, E ); \
    AN3 gate_BDF( BDF, B, D, F ); \
    AN3 gate_BEF( BEF, B, E, F ); \
    AN3 gate_CDE( CDE, C, D, E ); \
    AN3 gate_CDF( CDF, C, D, F ); \
    AN3 gate_CEF( CEF, C, E, F ); \
    AN3 gate_DEF( DEF, D, E, F );

`define wires_4_6 \
    wire  ABCD, ABCE, ABCF, ABDE, ABDF, ABEF, ACDE, ACDF, ACEF, ADEF, BCDE, BCDF, BCEF, BDEF, CDEF; \
    AN4 gate_ABCD( ABCD, A, B, C, D); \
    AN4 gate_ABCE( ABCE, A, B, C, E); \
    AN4 gate_ABCF( ABCF, A, B, C, F); \
    AN4 gate_ABDE( ABDE, A, B, D, E); \
    AN4 gate_ABDF( ABDF, A, B, D, F); \
    AN4 gate_ABEF( ABEF, A, B, E, F); \
    AN4 gate_ACDE( ACDE, A, C, D, E); \
    AN4 gate_ACDF( ACDF, A, C, D, F); \
    AN4 gate_ACEF( ACEF, A, C, E, F); \
    AN4 gate_ADEF( ADEF, A, D, E, F); \
    AN4 gate_BCDE( BCDE, B, C, D, E); \
    AN4 gate_BCDF( BCDF, B, C, D, F); \
    AN4 gate_BCEF( BCEF, B, C, E, F); \
    AN4 gate_BDEF( BDEF, B, D, E, F); \
    AN4 gate_CDEF( CDEF, C, D, E, F);

`define wires_5_6 \
    wire  BCDEF, ACDEF, ABDEF, ABCEF, ABCDF, ABCDE; \
    AN5 gate_BCDEF( BCDEF, B, C, D, E, F ); \
    AN5 gate_ACDEF( ACDEF, A, C, D, E, F ); \
    AN5 gate_ABDEF( ABDEF, A, B, D, E, F ); \
    AN5 gate_ABCEF( ABCEF, A, B, C, E, F ); \
    AN5 gate_ABCDF( ABCDF, A, B, C, D, F ); \
    AN5 gate_ABCDE( ABCDE, A, B, C, D, E );

`define wires_6_6 \
    wire  ABCDEF; \
    AN6 gate_ABCDEF( ABCDEF, A, B, C, D, E, F );

`define wires_2_5 \
    wire AB, AC, AD, AE, BC, BD, BE, CD, CE, DE; \
    AN2 gate_AB( AB, A, B ); \
    AN2 gate_AC( AC, A, C ); \
    AN2 gate_AD( AD, A, D ); \
    AN2 gate_AE( AE, A, E ); \
    AN2 gate_BC( BC, B, C ); \
    AN2 gate_BD( BD, B, D ); \
    AN2 gate_BE( BE, B, E ); \
    AN2 gate_CD( CD, C, D ); \
    AN2 gate_CE( CE, C, E ); \
    AN2 gate_DE( DE, D, E );

`define wires_3_5 \
    wire ABC, ABD, ABE, ACD, ACE, ADE, BCD, BCE, BDE, CDE; \
    AN3 gate_ABC( ABC, A, B, C); \
    AN3 gate_ABD( ABD, A, B, D); \
    AN3 gate_ABE( ABE, A, B, E); \
    AN3 gate_ACD( ACD, A, C, D); \
    AN3 gate_ACE( ACE, A, C, E); \
    AN3 gate_ADE( ADE, A, D, E); \
    AN3 gate_BCD( BCD, B, C, D); \
    AN3 gate_BCE( BCE, B, C, E); \
    AN3 gate_BDE( BDE, B, D, E); \
    AN3 gate_CDE( CDE, C, D, E);

`define wires_4_5 \
    wire BCDE, ACDE, ABDE, ABCE, ABCD; \
    AN4 gate_BCDE( BCDE, B, C, D, E); \
    AN4 gate_ACDE( ACDE, A, C, D, E); \
    AN4 gate_ABDE( ABDE, A, B, D, E); \
    AN4 gate_ABCE( ABCE, A, B, C, E); \
    AN4 gate_ABCD( ABCD, A, B, C, D);

`define wires_5_5 \
    wire ABCDE; \
    AN5 gate_ABCDE( ABCDE, A, B, C, D, E );

module Sanitizer( o, vec_63_bits);
    input  [62:0]   vec_63_bits;
    output [62:0]   o;
    wire   [1952:0] dummy;
    foobar f0( dummy[ 0], vec_63_bits[ 1], vec_63_bits[ 0] );
    foobar f1( dummy[ 1], vec_63_bits[ 2], vec_63_bits[ 0] );
    foobar f2( dummy[ 2], vec_63_bits[ 3], vec_63_bits[ 0] );
    foobar f3( dummy[ 3], vec_63_bits[ 4], vec_63_bits[ 0] );
    foobar f4( dummy[ 4], vec_63_bits[ 5], vec_63_bits[ 0] );
    foobar f5( dummy[ 5], vec_63_bits[ 6], vec_63_bits[ 0] );
    foobar f6( dummy[ 6], vec_63_bits[ 7], vec_63_bits[ 0] );
    foobar f7( dummy[ 7], vec_63_bits[ 8], vec_63_bits[ 0] );
    foobar f8( dummy[ 8], vec_63_bits[ 9], vec_63_bits[ 0] );
    foobar f9( dummy[ 9], vec_63_bits[10], vec_63_bits[ 0] );
    foobar f10( dummy[10], vec_63_bits[11], vec_63_bits[ 0] );
    foobar f11( dummy[11], vec_63_bits[12], vec_63_bits[ 0] );
    foobar f12( dummy[12], vec_63_bits[13], vec_63_bits[ 0] );
    foobar f13( dummy[13], vec_63_bits[14], vec_63_bits[ 0] );
    foobar f14( dummy[14], vec_63_bits[15], vec_63_bits[ 0] );
    foobar f15( dummy[15], vec_63_bits[16], vec_63_bits[ 0] );
    foobar f16( dummy[16], vec_63_bits[17], vec_63_bits[ 0] );
    foobar f17( dummy[17], vec_63_bits[18], vec_63_bits[ 0] );
    foobar f18( dummy[18], vec_63_bits[19], vec_63_bits[ 0] );
    foobar f19( dummy[19], vec_63_bits[20], vec_63_bits[ 0] );
    foobar f20( dummy[20], vec_63_bits[21], vec_63_bits[ 0] );
    foobar f21( dummy[21], vec_63_bits[22], vec_63_bits[ 0] );
    foobar f22( dummy[22], vec_63_bits[23], vec_63_bits[ 0] );
    foobar f23( dummy[23], vec_63_bits[24], vec_63_bits[ 0] );
    foobar f24( dummy[24], vec_63_bits[25], vec_63_bits[ 0] );
    foobar f25( dummy[25], vec_63_bits[26], vec_63_bits[ 0] );
    foobar f26( dummy[26], vec_63_bits[27], vec_63_bits[ 0] );
    foobar f27( dummy[27], vec_63_bits[28], vec_63_bits[ 0] );
    foobar f28( dummy[28], vec_63_bits[29], vec_63_bits[ 0] );
    foobar f29( dummy[29], vec_63_bits[30], vec_63_bits[ 0] );
    foobar f30( dummy[30], vec_63_bits[31], vec_63_bits[ 0] );
    foobar f31( dummy[31], vec_63_bits[32], vec_63_bits[ 0] );
    foobar f32( dummy[32], vec_63_bits[33], vec_63_bits[ 0] );
    foobar f33( dummy[33], vec_63_bits[34], vec_63_bits[ 0] );
    foobar f34( dummy[34], vec_63_bits[35], vec_63_bits[ 0] );
    foobar f35( dummy[35], vec_63_bits[36], vec_63_bits[ 0] );
    foobar f36( dummy[36], vec_63_bits[37], vec_63_bits[ 0] );
    foobar f37( dummy[37], vec_63_bits[38], vec_63_bits[ 0] );
    foobar f38( dummy[38], vec_63_bits[39], vec_63_bits[ 0] );
    foobar f39( dummy[39], vec_63_bits[40], vec_63_bits[ 0] );
    foobar f40( dummy[40], vec_63_bits[41], vec_63_bits[ 0] );
    foobar f41( dummy[41], vec_63_bits[42], vec_63_bits[ 0] );
    foobar f42( dummy[42], vec_63_bits[43], vec_63_bits[ 0] );
    foobar f43( dummy[43], vec_63_bits[44], vec_63_bits[ 0] );
    foobar f44( dummy[44], vec_63_bits[45], vec_63_bits[ 0] );
    foobar f45( dummy[45], vec_63_bits[46], vec_63_bits[ 0] );
    foobar f46( dummy[46], vec_63_bits[47], vec_63_bits[ 0] );
    foobar f47( dummy[47], vec_63_bits[48], vec_63_bits[ 0] );
    foobar f48( dummy[48], vec_63_bits[49], vec_63_bits[ 0] );
    foobar f49( dummy[49], vec_63_bits[50], vec_63_bits[ 0] );
    foobar f50( dummy[50], vec_63_bits[51], vec_63_bits[ 0] );
    foobar f51( dummy[51], vec_63_bits[52], vec_63_bits[ 0] );
    foobar f52( dummy[52], vec_63_bits[53], vec_63_bits[ 0] );
    foobar f53( dummy[53], vec_63_bits[54], vec_63_bits[ 0] );
    foobar f54( dummy[54], vec_63_bits[55], vec_63_bits[ 0] );
    foobar f55( dummy[55], vec_63_bits[56], vec_63_bits[ 0] );
    foobar f56( dummy[56], vec_63_bits[57], vec_63_bits[ 0] );
    foobar f57( dummy[57], vec_63_bits[58], vec_63_bits[ 0] );
    foobar f58( dummy[58], vec_63_bits[59], vec_63_bits[ 0] );
    foobar f59( dummy[59], vec_63_bits[60], vec_63_bits[ 0] );
    foobar f60( dummy[60], vec_63_bits[61], vec_63_bits[ 0] );
    foobar f61( dummy[61], vec_63_bits[62], vec_63_bits[ 0] );
    AN64   an0( o[0], {dummy[0], dummy[1], dummy[2], dummy[3], dummy[4], dummy[5], dummy[6], dummy[7], dummy[8], dummy[9], dummy[10], dummy[11], dummy[12], dummy[13], dummy[14], dummy[15], dummy[16], dummy[17], dummy[18], dummy[19], dummy[20], dummy[21], dummy[22], dummy[23], dummy[24], dummy[25], dummy[26], dummy[27], dummy[28], dummy[29], dummy[30], dummy[31], dummy[32], dummy[33], dummy[34], dummy[35], dummy[36], dummy[37], dummy[38], dummy[39], dummy[40], dummy[41], dummy[42], dummy[43], dummy[44], dummy[45], dummy[46], dummy[47], dummy[48], dummy[49], dummy[50], dummy[51], dummy[52], dummy[53], dummy[54], dummy[55], dummy[56], dummy[57], dummy[58], dummy[59], dummy[60], dummy[61], 1'b1, 1'b1 } );
    foobar f62( dummy[62], vec_63_bits[ 2], vec_63_bits[ 1] );
    foobar f63( dummy[63], vec_63_bits[ 3], vec_63_bits[ 1] );
    foobar f64( dummy[64], vec_63_bits[ 4], vec_63_bits[ 1] );
    foobar f65( dummy[65], vec_63_bits[ 5], vec_63_bits[ 1] );
    foobar f66( dummy[66], vec_63_bits[ 6], vec_63_bits[ 1] );
    foobar f67( dummy[67], vec_63_bits[ 7], vec_63_bits[ 1] );
    foobar f68( dummy[68], vec_63_bits[ 8], vec_63_bits[ 1] );
    foobar f69( dummy[69], vec_63_bits[ 9], vec_63_bits[ 1] );
    foobar f70( dummy[70], vec_63_bits[10], vec_63_bits[ 1] );
    foobar f71( dummy[71], vec_63_bits[11], vec_63_bits[ 1] );
    foobar f72( dummy[72], vec_63_bits[12], vec_63_bits[ 1] );
    foobar f73( dummy[73], vec_63_bits[13], vec_63_bits[ 1] );
    foobar f74( dummy[74], vec_63_bits[14], vec_63_bits[ 1] );
    foobar f75( dummy[75], vec_63_bits[15], vec_63_bits[ 1] );
    foobar f76( dummy[76], vec_63_bits[16], vec_63_bits[ 1] );
    foobar f77( dummy[77], vec_63_bits[17], vec_63_bits[ 1] );
    foobar f78( dummy[78], vec_63_bits[18], vec_63_bits[ 1] );
    foobar f79( dummy[79], vec_63_bits[19], vec_63_bits[ 1] );
    foobar f80( dummy[80], vec_63_bits[20], vec_63_bits[ 1] );
    foobar f81( dummy[81], vec_63_bits[21], vec_63_bits[ 1] );
    foobar f82( dummy[82], vec_63_bits[22], vec_63_bits[ 1] );
    foobar f83( dummy[83], vec_63_bits[23], vec_63_bits[ 1] );
    foobar f84( dummy[84], vec_63_bits[24], vec_63_bits[ 1] );
    foobar f85( dummy[85], vec_63_bits[25], vec_63_bits[ 1] );
    foobar f86( dummy[86], vec_63_bits[26], vec_63_bits[ 1] );
    foobar f87( dummy[87], vec_63_bits[27], vec_63_bits[ 1] );
    foobar f88( dummy[88], vec_63_bits[28], vec_63_bits[ 1] );
    foobar f89( dummy[89], vec_63_bits[29], vec_63_bits[ 1] );
    foobar f90( dummy[90], vec_63_bits[30], vec_63_bits[ 1] );
    foobar f91( dummy[91], vec_63_bits[31], vec_63_bits[ 1] );
    foobar f92( dummy[92], vec_63_bits[32], vec_63_bits[ 1] );
    foobar f93( dummy[93], vec_63_bits[33], vec_63_bits[ 1] );
    foobar f94( dummy[94], vec_63_bits[34], vec_63_bits[ 1] );
    foobar f95( dummy[95], vec_63_bits[35], vec_63_bits[ 1] );
    foobar f96( dummy[96], vec_63_bits[36], vec_63_bits[ 1] );
    foobar f97( dummy[97], vec_63_bits[37], vec_63_bits[ 1] );
    foobar f98( dummy[98], vec_63_bits[38], vec_63_bits[ 1] );
    foobar f99( dummy[99], vec_63_bits[39], vec_63_bits[ 1] );
    foobar f100( dummy[100], vec_63_bits[40], vec_63_bits[ 1] );
    foobar f101( dummy[101], vec_63_bits[41], vec_63_bits[ 1] );
    foobar f102( dummy[102], vec_63_bits[42], vec_63_bits[ 1] );
    foobar f103( dummy[103], vec_63_bits[43], vec_63_bits[ 1] );
    foobar f104( dummy[104], vec_63_bits[44], vec_63_bits[ 1] );
    foobar f105( dummy[105], vec_63_bits[45], vec_63_bits[ 1] );
    foobar f106( dummy[106], vec_63_bits[46], vec_63_bits[ 1] );
    foobar f107( dummy[107], vec_63_bits[47], vec_63_bits[ 1] );
    foobar f108( dummy[108], vec_63_bits[48], vec_63_bits[ 1] );
    foobar f109( dummy[109], vec_63_bits[49], vec_63_bits[ 1] );
    foobar f110( dummy[110], vec_63_bits[50], vec_63_bits[ 1] );
    foobar f111( dummy[111], vec_63_bits[51], vec_63_bits[ 1] );
    foobar f112( dummy[112], vec_63_bits[52], vec_63_bits[ 1] );
    foobar f113( dummy[113], vec_63_bits[53], vec_63_bits[ 1] );
    foobar f114( dummy[114], vec_63_bits[54], vec_63_bits[ 1] );
    foobar f115( dummy[115], vec_63_bits[55], vec_63_bits[ 1] );
    foobar f116( dummy[116], vec_63_bits[56], vec_63_bits[ 1] );
    foobar f117( dummy[117], vec_63_bits[57], vec_63_bits[ 1] );
    foobar f118( dummy[118], vec_63_bits[58], vec_63_bits[ 1] );
    foobar f119( dummy[119], vec_63_bits[59], vec_63_bits[ 1] );
    foobar f120( dummy[120], vec_63_bits[60], vec_63_bits[ 1] );
    foobar f121( dummy[121], vec_63_bits[61], vec_63_bits[ 1] );
    foobar f122( dummy[122], vec_63_bits[62], vec_63_bits[ 1] );
    AN64   an1( o[1], {dummy[62], dummy[63], dummy[64], dummy[65], dummy[66], dummy[67], dummy[68], dummy[69], dummy[70], dummy[71], dummy[72], dummy[73], dummy[74], dummy[75], dummy[76], dummy[77], dummy[78], dummy[79], dummy[80], dummy[81], dummy[82], dummy[83], dummy[84], dummy[85], dummy[86], dummy[87], dummy[88], dummy[89], dummy[90], dummy[91], dummy[92], dummy[93], dummy[94], dummy[95], dummy[96], dummy[97], dummy[98], dummy[99], dummy[100], dummy[101], dummy[102], dummy[103], dummy[104], dummy[105], dummy[106], dummy[107], dummy[108], dummy[109], dummy[110], dummy[111], dummy[112], dummy[113], dummy[114], dummy[115], dummy[116], dummy[117], dummy[118], dummy[119], dummy[120], dummy[121], dummy[122], 1'b1, 1'b1, 1'b1 } );
    foobar f123( dummy[123], vec_63_bits[ 3], vec_63_bits[ 2] );
    foobar f124( dummy[124], vec_63_bits[ 4], vec_63_bits[ 2] );
    foobar f125( dummy[125], vec_63_bits[ 5], vec_63_bits[ 2] );
    foobar f126( dummy[126], vec_63_bits[ 6], vec_63_bits[ 2] );
    foobar f127( dummy[127], vec_63_bits[ 7], vec_63_bits[ 2] );
    foobar f128( dummy[128], vec_63_bits[ 8], vec_63_bits[ 2] );
    foobar f129( dummy[129], vec_63_bits[ 9], vec_63_bits[ 2] );
    foobar f130( dummy[130], vec_63_bits[10], vec_63_bits[ 2] );
    foobar f131( dummy[131], vec_63_bits[11], vec_63_bits[ 2] );
    foobar f132( dummy[132], vec_63_bits[12], vec_63_bits[ 2] );
    foobar f133( dummy[133], vec_63_bits[13], vec_63_bits[ 2] );
    foobar f134( dummy[134], vec_63_bits[14], vec_63_bits[ 2] );
    foobar f135( dummy[135], vec_63_bits[15], vec_63_bits[ 2] );
    foobar f136( dummy[136], vec_63_bits[16], vec_63_bits[ 2] );
    foobar f137( dummy[137], vec_63_bits[17], vec_63_bits[ 2] );
    foobar f138( dummy[138], vec_63_bits[18], vec_63_bits[ 2] );
    foobar f139( dummy[139], vec_63_bits[19], vec_63_bits[ 2] );
    foobar f140( dummy[140], vec_63_bits[20], vec_63_bits[ 2] );
    foobar f141( dummy[141], vec_63_bits[21], vec_63_bits[ 2] );
    foobar f142( dummy[142], vec_63_bits[22], vec_63_bits[ 2] );
    foobar f143( dummy[143], vec_63_bits[23], vec_63_bits[ 2] );
    foobar f144( dummy[144], vec_63_bits[24], vec_63_bits[ 2] );
    foobar f145( dummy[145], vec_63_bits[25], vec_63_bits[ 2] );
    foobar f146( dummy[146], vec_63_bits[26], vec_63_bits[ 2] );
    foobar f147( dummy[147], vec_63_bits[27], vec_63_bits[ 2] );
    foobar f148( dummy[148], vec_63_bits[28], vec_63_bits[ 2] );
    foobar f149( dummy[149], vec_63_bits[29], vec_63_bits[ 2] );
    foobar f150( dummy[150], vec_63_bits[30], vec_63_bits[ 2] );
    foobar f151( dummy[151], vec_63_bits[31], vec_63_bits[ 2] );
    foobar f152( dummy[152], vec_63_bits[32], vec_63_bits[ 2] );
    foobar f153( dummy[153], vec_63_bits[33], vec_63_bits[ 2] );
    foobar f154( dummy[154], vec_63_bits[34], vec_63_bits[ 2] );
    foobar f155( dummy[155], vec_63_bits[35], vec_63_bits[ 2] );
    foobar f156( dummy[156], vec_63_bits[36], vec_63_bits[ 2] );
    foobar f157( dummy[157], vec_63_bits[37], vec_63_bits[ 2] );
    foobar f158( dummy[158], vec_63_bits[38], vec_63_bits[ 2] );
    foobar f159( dummy[159], vec_63_bits[39], vec_63_bits[ 2] );
    foobar f160( dummy[160], vec_63_bits[40], vec_63_bits[ 2] );
    foobar f161( dummy[161], vec_63_bits[41], vec_63_bits[ 2] );
    foobar f162( dummy[162], vec_63_bits[42], vec_63_bits[ 2] );
    foobar f163( dummy[163], vec_63_bits[43], vec_63_bits[ 2] );
    foobar f164( dummy[164], vec_63_bits[44], vec_63_bits[ 2] );
    foobar f165( dummy[165], vec_63_bits[45], vec_63_bits[ 2] );
    foobar f166( dummy[166], vec_63_bits[46], vec_63_bits[ 2] );
    foobar f167( dummy[167], vec_63_bits[47], vec_63_bits[ 2] );
    foobar f168( dummy[168], vec_63_bits[48], vec_63_bits[ 2] );
    foobar f169( dummy[169], vec_63_bits[49], vec_63_bits[ 2] );
    foobar f170( dummy[170], vec_63_bits[50], vec_63_bits[ 2] );
    foobar f171( dummy[171], vec_63_bits[51], vec_63_bits[ 2] );
    foobar f172( dummy[172], vec_63_bits[52], vec_63_bits[ 2] );
    foobar f173( dummy[173], vec_63_bits[53], vec_63_bits[ 2] );
    foobar f174( dummy[174], vec_63_bits[54], vec_63_bits[ 2] );
    foobar f175( dummy[175], vec_63_bits[55], vec_63_bits[ 2] );
    foobar f176( dummy[176], vec_63_bits[56], vec_63_bits[ 2] );
    foobar f177( dummy[177], vec_63_bits[57], vec_63_bits[ 2] );
    foobar f178( dummy[178], vec_63_bits[58], vec_63_bits[ 2] );
    foobar f179( dummy[179], vec_63_bits[59], vec_63_bits[ 2] );
    foobar f180( dummy[180], vec_63_bits[60], vec_63_bits[ 2] );
    foobar f181( dummy[181], vec_63_bits[61], vec_63_bits[ 2] );
    foobar f182( dummy[182], vec_63_bits[62], vec_63_bits[ 2] );
    AN64   an2( o[2], {dummy[123], dummy[124], dummy[125], dummy[126], dummy[127], dummy[128], dummy[129], dummy[130], dummy[131], dummy[132], dummy[133], dummy[134], dummy[135], dummy[136], dummy[137], dummy[138], dummy[139], dummy[140], dummy[141], dummy[142], dummy[143], dummy[144], dummy[145], dummy[146], dummy[147], dummy[148], dummy[149], dummy[150], dummy[151], dummy[152], dummy[153], dummy[154], dummy[155], dummy[156], dummy[157], dummy[158], dummy[159], dummy[160], dummy[161], dummy[162], dummy[163], dummy[164], dummy[165], dummy[166], dummy[167], dummy[168], dummy[169], dummy[170], dummy[171], dummy[172], dummy[173], dummy[174], dummy[175], dummy[176], dummy[177], dummy[178], dummy[179], dummy[180], dummy[181], dummy[182], 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f183( dummy[183], vec_63_bits[ 4], vec_63_bits[ 3] );
    foobar f184( dummy[184], vec_63_bits[ 5], vec_63_bits[ 3] );
    foobar f185( dummy[185], vec_63_bits[ 6], vec_63_bits[ 3] );
    foobar f186( dummy[186], vec_63_bits[ 7], vec_63_bits[ 3] );
    foobar f187( dummy[187], vec_63_bits[ 8], vec_63_bits[ 3] );
    foobar f188( dummy[188], vec_63_bits[ 9], vec_63_bits[ 3] );
    foobar f189( dummy[189], vec_63_bits[10], vec_63_bits[ 3] );
    foobar f190( dummy[190], vec_63_bits[11], vec_63_bits[ 3] );
    foobar f191( dummy[191], vec_63_bits[12], vec_63_bits[ 3] );
    foobar f192( dummy[192], vec_63_bits[13], vec_63_bits[ 3] );
    foobar f193( dummy[193], vec_63_bits[14], vec_63_bits[ 3] );
    foobar f194( dummy[194], vec_63_bits[15], vec_63_bits[ 3] );
    foobar f195( dummy[195], vec_63_bits[16], vec_63_bits[ 3] );
    foobar f196( dummy[196], vec_63_bits[17], vec_63_bits[ 3] );
    foobar f197( dummy[197], vec_63_bits[18], vec_63_bits[ 3] );
    foobar f198( dummy[198], vec_63_bits[19], vec_63_bits[ 3] );
    foobar f199( dummy[199], vec_63_bits[20], vec_63_bits[ 3] );
    foobar f200( dummy[200], vec_63_bits[21], vec_63_bits[ 3] );
    foobar f201( dummy[201], vec_63_bits[22], vec_63_bits[ 3] );
    foobar f202( dummy[202], vec_63_bits[23], vec_63_bits[ 3] );
    foobar f203( dummy[203], vec_63_bits[24], vec_63_bits[ 3] );
    foobar f204( dummy[204], vec_63_bits[25], vec_63_bits[ 3] );
    foobar f205( dummy[205], vec_63_bits[26], vec_63_bits[ 3] );
    foobar f206( dummy[206], vec_63_bits[27], vec_63_bits[ 3] );
    foobar f207( dummy[207], vec_63_bits[28], vec_63_bits[ 3] );
    foobar f208( dummy[208], vec_63_bits[29], vec_63_bits[ 3] );
    foobar f209( dummy[209], vec_63_bits[30], vec_63_bits[ 3] );
    foobar f210( dummy[210], vec_63_bits[31], vec_63_bits[ 3] );
    foobar f211( dummy[211], vec_63_bits[32], vec_63_bits[ 3] );
    foobar f212( dummy[212], vec_63_bits[33], vec_63_bits[ 3] );
    foobar f213( dummy[213], vec_63_bits[34], vec_63_bits[ 3] );
    foobar f214( dummy[214], vec_63_bits[35], vec_63_bits[ 3] );
    foobar f215( dummy[215], vec_63_bits[36], vec_63_bits[ 3] );
    foobar f216( dummy[216], vec_63_bits[37], vec_63_bits[ 3] );
    foobar f217( dummy[217], vec_63_bits[38], vec_63_bits[ 3] );
    foobar f218( dummy[218], vec_63_bits[39], vec_63_bits[ 3] );
    foobar f219( dummy[219], vec_63_bits[40], vec_63_bits[ 3] );
    foobar f220( dummy[220], vec_63_bits[41], vec_63_bits[ 3] );
    foobar f221( dummy[221], vec_63_bits[42], vec_63_bits[ 3] );
    foobar f222( dummy[222], vec_63_bits[43], vec_63_bits[ 3] );
    foobar f223( dummy[223], vec_63_bits[44], vec_63_bits[ 3] );
    foobar f224( dummy[224], vec_63_bits[45], vec_63_bits[ 3] );
    foobar f225( dummy[225], vec_63_bits[46], vec_63_bits[ 3] );
    foobar f226( dummy[226], vec_63_bits[47], vec_63_bits[ 3] );
    foobar f227( dummy[227], vec_63_bits[48], vec_63_bits[ 3] );
    foobar f228( dummy[228], vec_63_bits[49], vec_63_bits[ 3] );
    foobar f229( dummy[229], vec_63_bits[50], vec_63_bits[ 3] );
    foobar f230( dummy[230], vec_63_bits[51], vec_63_bits[ 3] );
    foobar f231( dummy[231], vec_63_bits[52], vec_63_bits[ 3] );
    foobar f232( dummy[232], vec_63_bits[53], vec_63_bits[ 3] );
    foobar f233( dummy[233], vec_63_bits[54], vec_63_bits[ 3] );
    foobar f234( dummy[234], vec_63_bits[55], vec_63_bits[ 3] );
    foobar f235( dummy[235], vec_63_bits[56], vec_63_bits[ 3] );
    foobar f236( dummy[236], vec_63_bits[57], vec_63_bits[ 3] );
    foobar f237( dummy[237], vec_63_bits[58], vec_63_bits[ 3] );
    foobar f238( dummy[238], vec_63_bits[59], vec_63_bits[ 3] );
    foobar f239( dummy[239], vec_63_bits[60], vec_63_bits[ 3] );
    foobar f240( dummy[240], vec_63_bits[61], vec_63_bits[ 3] );
    foobar f241( dummy[241], vec_63_bits[62], vec_63_bits[ 3] );
    AN64   an3( o[3], {dummy[183], dummy[184], dummy[185], dummy[186], dummy[187], dummy[188], dummy[189], dummy[190], dummy[191], dummy[192], dummy[193], dummy[194], dummy[195], dummy[196], dummy[197], dummy[198], dummy[199], dummy[200], dummy[201], dummy[202], dummy[203], dummy[204], dummy[205], dummy[206], dummy[207], dummy[208], dummy[209], dummy[210], dummy[211], dummy[212], dummy[213], dummy[214], dummy[215], dummy[216], dummy[217], dummy[218], dummy[219], dummy[220], dummy[221], dummy[222], dummy[223], dummy[224], dummy[225], dummy[226], dummy[227], dummy[228], dummy[229], dummy[230], dummy[231], dummy[232], dummy[233], dummy[234], dummy[235], dummy[236], dummy[237], dummy[238], dummy[239], dummy[240], dummy[241], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f242( dummy[242], vec_63_bits[ 5], vec_63_bits[ 4] );
    foobar f243( dummy[243], vec_63_bits[ 6], vec_63_bits[ 4] );
    foobar f244( dummy[244], vec_63_bits[ 7], vec_63_bits[ 4] );
    foobar f245( dummy[245], vec_63_bits[ 8], vec_63_bits[ 4] );
    foobar f246( dummy[246], vec_63_bits[ 9], vec_63_bits[ 4] );
    foobar f247( dummy[247], vec_63_bits[10], vec_63_bits[ 4] );
    foobar f248( dummy[248], vec_63_bits[11], vec_63_bits[ 4] );
    foobar f249( dummy[249], vec_63_bits[12], vec_63_bits[ 4] );
    foobar f250( dummy[250], vec_63_bits[13], vec_63_bits[ 4] );
    foobar f251( dummy[251], vec_63_bits[14], vec_63_bits[ 4] );
    foobar f252( dummy[252], vec_63_bits[15], vec_63_bits[ 4] );
    foobar f253( dummy[253], vec_63_bits[16], vec_63_bits[ 4] );
    foobar f254( dummy[254], vec_63_bits[17], vec_63_bits[ 4] );
    foobar f255( dummy[255], vec_63_bits[18], vec_63_bits[ 4] );
    foobar f256( dummy[256], vec_63_bits[19], vec_63_bits[ 4] );
    foobar f257( dummy[257], vec_63_bits[20], vec_63_bits[ 4] );
    foobar f258( dummy[258], vec_63_bits[21], vec_63_bits[ 4] );
    foobar f259( dummy[259], vec_63_bits[22], vec_63_bits[ 4] );
    foobar f260( dummy[260], vec_63_bits[23], vec_63_bits[ 4] );
    foobar f261( dummy[261], vec_63_bits[24], vec_63_bits[ 4] );
    foobar f262( dummy[262], vec_63_bits[25], vec_63_bits[ 4] );
    foobar f263( dummy[263], vec_63_bits[26], vec_63_bits[ 4] );
    foobar f264( dummy[264], vec_63_bits[27], vec_63_bits[ 4] );
    foobar f265( dummy[265], vec_63_bits[28], vec_63_bits[ 4] );
    foobar f266( dummy[266], vec_63_bits[29], vec_63_bits[ 4] );
    foobar f267( dummy[267], vec_63_bits[30], vec_63_bits[ 4] );
    foobar f268( dummy[268], vec_63_bits[31], vec_63_bits[ 4] );
    foobar f269( dummy[269], vec_63_bits[32], vec_63_bits[ 4] );
    foobar f270( dummy[270], vec_63_bits[33], vec_63_bits[ 4] );
    foobar f271( dummy[271], vec_63_bits[34], vec_63_bits[ 4] );
    foobar f272( dummy[272], vec_63_bits[35], vec_63_bits[ 4] );
    foobar f273( dummy[273], vec_63_bits[36], vec_63_bits[ 4] );
    foobar f274( dummy[274], vec_63_bits[37], vec_63_bits[ 4] );
    foobar f275( dummy[275], vec_63_bits[38], vec_63_bits[ 4] );
    foobar f276( dummy[276], vec_63_bits[39], vec_63_bits[ 4] );
    foobar f277( dummy[277], vec_63_bits[40], vec_63_bits[ 4] );
    foobar f278( dummy[278], vec_63_bits[41], vec_63_bits[ 4] );
    foobar f279( dummy[279], vec_63_bits[42], vec_63_bits[ 4] );
    foobar f280( dummy[280], vec_63_bits[43], vec_63_bits[ 4] );
    foobar f281( dummy[281], vec_63_bits[44], vec_63_bits[ 4] );
    foobar f282( dummy[282], vec_63_bits[45], vec_63_bits[ 4] );
    foobar f283( dummy[283], vec_63_bits[46], vec_63_bits[ 4] );
    foobar f284( dummy[284], vec_63_bits[47], vec_63_bits[ 4] );
    foobar f285( dummy[285], vec_63_bits[48], vec_63_bits[ 4] );
    foobar f286( dummy[286], vec_63_bits[49], vec_63_bits[ 4] );
    foobar f287( dummy[287], vec_63_bits[50], vec_63_bits[ 4] );
    foobar f288( dummy[288], vec_63_bits[51], vec_63_bits[ 4] );
    foobar f289( dummy[289], vec_63_bits[52], vec_63_bits[ 4] );
    foobar f290( dummy[290], vec_63_bits[53], vec_63_bits[ 4] );
    foobar f291( dummy[291], vec_63_bits[54], vec_63_bits[ 4] );
    foobar f292( dummy[292], vec_63_bits[55], vec_63_bits[ 4] );
    foobar f293( dummy[293], vec_63_bits[56], vec_63_bits[ 4] );
    foobar f294( dummy[294], vec_63_bits[57], vec_63_bits[ 4] );
    foobar f295( dummy[295], vec_63_bits[58], vec_63_bits[ 4] );
    foobar f296( dummy[296], vec_63_bits[59], vec_63_bits[ 4] );
    foobar f297( dummy[297], vec_63_bits[60], vec_63_bits[ 4] );
    foobar f298( dummy[298], vec_63_bits[61], vec_63_bits[ 4] );
    foobar f299( dummy[299], vec_63_bits[62], vec_63_bits[ 4] );
    AN64   an4( o[4], {dummy[242], dummy[243], dummy[244], dummy[245], dummy[246], dummy[247], dummy[248], dummy[249], dummy[250], dummy[251], dummy[252], dummy[253], dummy[254], dummy[255], dummy[256], dummy[257], dummy[258], dummy[259], dummy[260], dummy[261], dummy[262], dummy[263], dummy[264], dummy[265], dummy[266], dummy[267], dummy[268], dummy[269], dummy[270], dummy[271], dummy[272], dummy[273], dummy[274], dummy[275], dummy[276], dummy[277], dummy[278], dummy[279], dummy[280], dummy[281], dummy[282], dummy[283], dummy[284], dummy[285], dummy[286], dummy[287], dummy[288], dummy[289], dummy[290], dummy[291], dummy[292], dummy[293], dummy[294], dummy[295], dummy[296], dummy[297], dummy[298], dummy[299], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f300( dummy[300], vec_63_bits[ 6], vec_63_bits[ 5] );
    foobar f301( dummy[301], vec_63_bits[ 7], vec_63_bits[ 5] );
    foobar f302( dummy[302], vec_63_bits[ 8], vec_63_bits[ 5] );
    foobar f303( dummy[303], vec_63_bits[ 9], vec_63_bits[ 5] );
    foobar f304( dummy[304], vec_63_bits[10], vec_63_bits[ 5] );
    foobar f305( dummy[305], vec_63_bits[11], vec_63_bits[ 5] );
    foobar f306( dummy[306], vec_63_bits[12], vec_63_bits[ 5] );
    foobar f307( dummy[307], vec_63_bits[13], vec_63_bits[ 5] );
    foobar f308( dummy[308], vec_63_bits[14], vec_63_bits[ 5] );
    foobar f309( dummy[309], vec_63_bits[15], vec_63_bits[ 5] );
    foobar f310( dummy[310], vec_63_bits[16], vec_63_bits[ 5] );
    foobar f311( dummy[311], vec_63_bits[17], vec_63_bits[ 5] );
    foobar f312( dummy[312], vec_63_bits[18], vec_63_bits[ 5] );
    foobar f313( dummy[313], vec_63_bits[19], vec_63_bits[ 5] );
    foobar f314( dummy[314], vec_63_bits[20], vec_63_bits[ 5] );
    foobar f315( dummy[315], vec_63_bits[21], vec_63_bits[ 5] );
    foobar f316( dummy[316], vec_63_bits[22], vec_63_bits[ 5] );
    foobar f317( dummy[317], vec_63_bits[23], vec_63_bits[ 5] );
    foobar f318( dummy[318], vec_63_bits[24], vec_63_bits[ 5] );
    foobar f319( dummy[319], vec_63_bits[25], vec_63_bits[ 5] );
    foobar f320( dummy[320], vec_63_bits[26], vec_63_bits[ 5] );
    foobar f321( dummy[321], vec_63_bits[27], vec_63_bits[ 5] );
    foobar f322( dummy[322], vec_63_bits[28], vec_63_bits[ 5] );
    foobar f323( dummy[323], vec_63_bits[29], vec_63_bits[ 5] );
    foobar f324( dummy[324], vec_63_bits[30], vec_63_bits[ 5] );
    foobar f325( dummy[325], vec_63_bits[31], vec_63_bits[ 5] );
    foobar f326( dummy[326], vec_63_bits[32], vec_63_bits[ 5] );
    foobar f327( dummy[327], vec_63_bits[33], vec_63_bits[ 5] );
    foobar f328( dummy[328], vec_63_bits[34], vec_63_bits[ 5] );
    foobar f329( dummy[329], vec_63_bits[35], vec_63_bits[ 5] );
    foobar f330( dummy[330], vec_63_bits[36], vec_63_bits[ 5] );
    foobar f331( dummy[331], vec_63_bits[37], vec_63_bits[ 5] );
    foobar f332( dummy[332], vec_63_bits[38], vec_63_bits[ 5] );
    foobar f333( dummy[333], vec_63_bits[39], vec_63_bits[ 5] );
    foobar f334( dummy[334], vec_63_bits[40], vec_63_bits[ 5] );
    foobar f335( dummy[335], vec_63_bits[41], vec_63_bits[ 5] );
    foobar f336( dummy[336], vec_63_bits[42], vec_63_bits[ 5] );
    foobar f337( dummy[337], vec_63_bits[43], vec_63_bits[ 5] );
    foobar f338( dummy[338], vec_63_bits[44], vec_63_bits[ 5] );
    foobar f339( dummy[339], vec_63_bits[45], vec_63_bits[ 5] );
    foobar f340( dummy[340], vec_63_bits[46], vec_63_bits[ 5] );
    foobar f341( dummy[341], vec_63_bits[47], vec_63_bits[ 5] );
    foobar f342( dummy[342], vec_63_bits[48], vec_63_bits[ 5] );
    foobar f343( dummy[343], vec_63_bits[49], vec_63_bits[ 5] );
    foobar f344( dummy[344], vec_63_bits[50], vec_63_bits[ 5] );
    foobar f345( dummy[345], vec_63_bits[51], vec_63_bits[ 5] );
    foobar f346( dummy[346], vec_63_bits[52], vec_63_bits[ 5] );
    foobar f347( dummy[347], vec_63_bits[53], vec_63_bits[ 5] );
    foobar f348( dummy[348], vec_63_bits[54], vec_63_bits[ 5] );
    foobar f349( dummy[349], vec_63_bits[55], vec_63_bits[ 5] );
    foobar f350( dummy[350], vec_63_bits[56], vec_63_bits[ 5] );
    foobar f351( dummy[351], vec_63_bits[57], vec_63_bits[ 5] );
    foobar f352( dummy[352], vec_63_bits[58], vec_63_bits[ 5] );
    foobar f353( dummy[353], vec_63_bits[59], vec_63_bits[ 5] );
    foobar f354( dummy[354], vec_63_bits[60], vec_63_bits[ 5] );
    foobar f355( dummy[355], vec_63_bits[61], vec_63_bits[ 5] );
    foobar f356( dummy[356], vec_63_bits[62], vec_63_bits[ 5] );
    AN64   an5( o[5], {dummy[300], dummy[301], dummy[302], dummy[303], dummy[304], dummy[305], dummy[306], dummy[307], dummy[308], dummy[309], dummy[310], dummy[311], dummy[312], dummy[313], dummy[314], dummy[315], dummy[316], dummy[317], dummy[318], dummy[319], dummy[320], dummy[321], dummy[322], dummy[323], dummy[324], dummy[325], dummy[326], dummy[327], dummy[328], dummy[329], dummy[330], dummy[331], dummy[332], dummy[333], dummy[334], dummy[335], dummy[336], dummy[337], dummy[338], dummy[339], dummy[340], dummy[341], dummy[342], dummy[343], dummy[344], dummy[345], dummy[346], dummy[347], dummy[348], dummy[349], dummy[350], dummy[351], dummy[352], dummy[353], dummy[354], dummy[355], dummy[356], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f357( dummy[357], vec_63_bits[ 7], vec_63_bits[ 6] );
    foobar f358( dummy[358], vec_63_bits[ 8], vec_63_bits[ 6] );
    foobar f359( dummy[359], vec_63_bits[ 9], vec_63_bits[ 6] );
    foobar f360( dummy[360], vec_63_bits[10], vec_63_bits[ 6] );
    foobar f361( dummy[361], vec_63_bits[11], vec_63_bits[ 6] );
    foobar f362( dummy[362], vec_63_bits[12], vec_63_bits[ 6] );
    foobar f363( dummy[363], vec_63_bits[13], vec_63_bits[ 6] );
    foobar f364( dummy[364], vec_63_bits[14], vec_63_bits[ 6] );
    foobar f365( dummy[365], vec_63_bits[15], vec_63_bits[ 6] );
    foobar f366( dummy[366], vec_63_bits[16], vec_63_bits[ 6] );
    foobar f367( dummy[367], vec_63_bits[17], vec_63_bits[ 6] );
    foobar f368( dummy[368], vec_63_bits[18], vec_63_bits[ 6] );
    foobar f369( dummy[369], vec_63_bits[19], vec_63_bits[ 6] );
    foobar f370( dummy[370], vec_63_bits[20], vec_63_bits[ 6] );
    foobar f371( dummy[371], vec_63_bits[21], vec_63_bits[ 6] );
    foobar f372( dummy[372], vec_63_bits[22], vec_63_bits[ 6] );
    foobar f373( dummy[373], vec_63_bits[23], vec_63_bits[ 6] );
    foobar f374( dummy[374], vec_63_bits[24], vec_63_bits[ 6] );
    foobar f375( dummy[375], vec_63_bits[25], vec_63_bits[ 6] );
    foobar f376( dummy[376], vec_63_bits[26], vec_63_bits[ 6] );
    foobar f377( dummy[377], vec_63_bits[27], vec_63_bits[ 6] );
    foobar f378( dummy[378], vec_63_bits[28], vec_63_bits[ 6] );
    foobar f379( dummy[379], vec_63_bits[29], vec_63_bits[ 6] );
    foobar f380( dummy[380], vec_63_bits[30], vec_63_bits[ 6] );
    foobar f381( dummy[381], vec_63_bits[31], vec_63_bits[ 6] );
    foobar f382( dummy[382], vec_63_bits[32], vec_63_bits[ 6] );
    foobar f383( dummy[383], vec_63_bits[33], vec_63_bits[ 6] );
    foobar f384( dummy[384], vec_63_bits[34], vec_63_bits[ 6] );
    foobar f385( dummy[385], vec_63_bits[35], vec_63_bits[ 6] );
    foobar f386( dummy[386], vec_63_bits[36], vec_63_bits[ 6] );
    foobar f387( dummy[387], vec_63_bits[37], vec_63_bits[ 6] );
    foobar f388( dummy[388], vec_63_bits[38], vec_63_bits[ 6] );
    foobar f389( dummy[389], vec_63_bits[39], vec_63_bits[ 6] );
    foobar f390( dummy[390], vec_63_bits[40], vec_63_bits[ 6] );
    foobar f391( dummy[391], vec_63_bits[41], vec_63_bits[ 6] );
    foobar f392( dummy[392], vec_63_bits[42], vec_63_bits[ 6] );
    foobar f393( dummy[393], vec_63_bits[43], vec_63_bits[ 6] );
    foobar f394( dummy[394], vec_63_bits[44], vec_63_bits[ 6] );
    foobar f395( dummy[395], vec_63_bits[45], vec_63_bits[ 6] );
    foobar f396( dummy[396], vec_63_bits[46], vec_63_bits[ 6] );
    foobar f397( dummy[397], vec_63_bits[47], vec_63_bits[ 6] );
    foobar f398( dummy[398], vec_63_bits[48], vec_63_bits[ 6] );
    foobar f399( dummy[399], vec_63_bits[49], vec_63_bits[ 6] );
    foobar f400( dummy[400], vec_63_bits[50], vec_63_bits[ 6] );
    foobar f401( dummy[401], vec_63_bits[51], vec_63_bits[ 6] );
    foobar f402( dummy[402], vec_63_bits[52], vec_63_bits[ 6] );
    foobar f403( dummy[403], vec_63_bits[53], vec_63_bits[ 6] );
    foobar f404( dummy[404], vec_63_bits[54], vec_63_bits[ 6] );
    foobar f405( dummy[405], vec_63_bits[55], vec_63_bits[ 6] );
    foobar f406( dummy[406], vec_63_bits[56], vec_63_bits[ 6] );
    foobar f407( dummy[407], vec_63_bits[57], vec_63_bits[ 6] );
    foobar f408( dummy[408], vec_63_bits[58], vec_63_bits[ 6] );
    foobar f409( dummy[409], vec_63_bits[59], vec_63_bits[ 6] );
    foobar f410( dummy[410], vec_63_bits[60], vec_63_bits[ 6] );
    foobar f411( dummy[411], vec_63_bits[61], vec_63_bits[ 6] );
    foobar f412( dummy[412], vec_63_bits[62], vec_63_bits[ 6] );
    AN64   an6( o[6], {dummy[357], dummy[358], dummy[359], dummy[360], dummy[361], dummy[362], dummy[363], dummy[364], dummy[365], dummy[366], dummy[367], dummy[368], dummy[369], dummy[370], dummy[371], dummy[372], dummy[373], dummy[374], dummy[375], dummy[376], dummy[377], dummy[378], dummy[379], dummy[380], dummy[381], dummy[382], dummy[383], dummy[384], dummy[385], dummy[386], dummy[387], dummy[388], dummy[389], dummy[390], dummy[391], dummy[392], dummy[393], dummy[394], dummy[395], dummy[396], dummy[397], dummy[398], dummy[399], dummy[400], dummy[401], dummy[402], dummy[403], dummy[404], dummy[405], dummy[406], dummy[407], dummy[408], dummy[409], dummy[410], dummy[411], dummy[412], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f413( dummy[413], vec_63_bits[ 8], vec_63_bits[ 7] );
    foobar f414( dummy[414], vec_63_bits[ 9], vec_63_bits[ 7] );
    foobar f415( dummy[415], vec_63_bits[10], vec_63_bits[ 7] );
    foobar f416( dummy[416], vec_63_bits[11], vec_63_bits[ 7] );
    foobar f417( dummy[417], vec_63_bits[12], vec_63_bits[ 7] );
    foobar f418( dummy[418], vec_63_bits[13], vec_63_bits[ 7] );
    foobar f419( dummy[419], vec_63_bits[14], vec_63_bits[ 7] );
    foobar f420( dummy[420], vec_63_bits[15], vec_63_bits[ 7] );
    foobar f421( dummy[421], vec_63_bits[16], vec_63_bits[ 7] );
    foobar f422( dummy[422], vec_63_bits[17], vec_63_bits[ 7] );
    foobar f423( dummy[423], vec_63_bits[18], vec_63_bits[ 7] );
    foobar f424( dummy[424], vec_63_bits[19], vec_63_bits[ 7] );
    foobar f425( dummy[425], vec_63_bits[20], vec_63_bits[ 7] );
    foobar f426( dummy[426], vec_63_bits[21], vec_63_bits[ 7] );
    foobar f427( dummy[427], vec_63_bits[22], vec_63_bits[ 7] );
    foobar f428( dummy[428], vec_63_bits[23], vec_63_bits[ 7] );
    foobar f429( dummy[429], vec_63_bits[24], vec_63_bits[ 7] );
    foobar f430( dummy[430], vec_63_bits[25], vec_63_bits[ 7] );
    foobar f431( dummy[431], vec_63_bits[26], vec_63_bits[ 7] );
    foobar f432( dummy[432], vec_63_bits[27], vec_63_bits[ 7] );
    foobar f433( dummy[433], vec_63_bits[28], vec_63_bits[ 7] );
    foobar f434( dummy[434], vec_63_bits[29], vec_63_bits[ 7] );
    foobar f435( dummy[435], vec_63_bits[30], vec_63_bits[ 7] );
    foobar f436( dummy[436], vec_63_bits[31], vec_63_bits[ 7] );
    foobar f437( dummy[437], vec_63_bits[32], vec_63_bits[ 7] );
    foobar f438( dummy[438], vec_63_bits[33], vec_63_bits[ 7] );
    foobar f439( dummy[439], vec_63_bits[34], vec_63_bits[ 7] );
    foobar f440( dummy[440], vec_63_bits[35], vec_63_bits[ 7] );
    foobar f441( dummy[441], vec_63_bits[36], vec_63_bits[ 7] );
    foobar f442( dummy[442], vec_63_bits[37], vec_63_bits[ 7] );
    foobar f443( dummy[443], vec_63_bits[38], vec_63_bits[ 7] );
    foobar f444( dummy[444], vec_63_bits[39], vec_63_bits[ 7] );
    foobar f445( dummy[445], vec_63_bits[40], vec_63_bits[ 7] );
    foobar f446( dummy[446], vec_63_bits[41], vec_63_bits[ 7] );
    foobar f447( dummy[447], vec_63_bits[42], vec_63_bits[ 7] );
    foobar f448( dummy[448], vec_63_bits[43], vec_63_bits[ 7] );
    foobar f449( dummy[449], vec_63_bits[44], vec_63_bits[ 7] );
    foobar f450( dummy[450], vec_63_bits[45], vec_63_bits[ 7] );
    foobar f451( dummy[451], vec_63_bits[46], vec_63_bits[ 7] );
    foobar f452( dummy[452], vec_63_bits[47], vec_63_bits[ 7] );
    foobar f453( dummy[453], vec_63_bits[48], vec_63_bits[ 7] );
    foobar f454( dummy[454], vec_63_bits[49], vec_63_bits[ 7] );
    foobar f455( dummy[455], vec_63_bits[50], vec_63_bits[ 7] );
    foobar f456( dummy[456], vec_63_bits[51], vec_63_bits[ 7] );
    foobar f457( dummy[457], vec_63_bits[52], vec_63_bits[ 7] );
    foobar f458( dummy[458], vec_63_bits[53], vec_63_bits[ 7] );
    foobar f459( dummy[459], vec_63_bits[54], vec_63_bits[ 7] );
    foobar f460( dummy[460], vec_63_bits[55], vec_63_bits[ 7] );
    foobar f461( dummy[461], vec_63_bits[56], vec_63_bits[ 7] );
    foobar f462( dummy[462], vec_63_bits[57], vec_63_bits[ 7] );
    foobar f463( dummy[463], vec_63_bits[58], vec_63_bits[ 7] );
    foobar f464( dummy[464], vec_63_bits[59], vec_63_bits[ 7] );
    foobar f465( dummy[465], vec_63_bits[60], vec_63_bits[ 7] );
    foobar f466( dummy[466], vec_63_bits[61], vec_63_bits[ 7] );
    foobar f467( dummy[467], vec_63_bits[62], vec_63_bits[ 7] );
    AN64   an7( o[7], {dummy[413], dummy[414], dummy[415], dummy[416], dummy[417], dummy[418], dummy[419], dummy[420], dummy[421], dummy[422], dummy[423], dummy[424], dummy[425], dummy[426], dummy[427], dummy[428], dummy[429], dummy[430], dummy[431], dummy[432], dummy[433], dummy[434], dummy[435], dummy[436], dummy[437], dummy[438], dummy[439], dummy[440], dummy[441], dummy[442], dummy[443], dummy[444], dummy[445], dummy[446], dummy[447], dummy[448], dummy[449], dummy[450], dummy[451], dummy[452], dummy[453], dummy[454], dummy[455], dummy[456], dummy[457], dummy[458], dummy[459], dummy[460], dummy[461], dummy[462], dummy[463], dummy[464], dummy[465], dummy[466], dummy[467], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f468( dummy[468], vec_63_bits[ 9], vec_63_bits[ 8] );
    foobar f469( dummy[469], vec_63_bits[10], vec_63_bits[ 8] );
    foobar f470( dummy[470], vec_63_bits[11], vec_63_bits[ 8] );
    foobar f471( dummy[471], vec_63_bits[12], vec_63_bits[ 8] );
    foobar f472( dummy[472], vec_63_bits[13], vec_63_bits[ 8] );
    foobar f473( dummy[473], vec_63_bits[14], vec_63_bits[ 8] );
    foobar f474( dummy[474], vec_63_bits[15], vec_63_bits[ 8] );
    foobar f475( dummy[475], vec_63_bits[16], vec_63_bits[ 8] );
    foobar f476( dummy[476], vec_63_bits[17], vec_63_bits[ 8] );
    foobar f477( dummy[477], vec_63_bits[18], vec_63_bits[ 8] );
    foobar f478( dummy[478], vec_63_bits[19], vec_63_bits[ 8] );
    foobar f479( dummy[479], vec_63_bits[20], vec_63_bits[ 8] );
    foobar f480( dummy[480], vec_63_bits[21], vec_63_bits[ 8] );
    foobar f481( dummy[481], vec_63_bits[22], vec_63_bits[ 8] );
    foobar f482( dummy[482], vec_63_bits[23], vec_63_bits[ 8] );
    foobar f483( dummy[483], vec_63_bits[24], vec_63_bits[ 8] );
    foobar f484( dummy[484], vec_63_bits[25], vec_63_bits[ 8] );
    foobar f485( dummy[485], vec_63_bits[26], vec_63_bits[ 8] );
    foobar f486( dummy[486], vec_63_bits[27], vec_63_bits[ 8] );
    foobar f487( dummy[487], vec_63_bits[28], vec_63_bits[ 8] );
    foobar f488( dummy[488], vec_63_bits[29], vec_63_bits[ 8] );
    foobar f489( dummy[489], vec_63_bits[30], vec_63_bits[ 8] );
    foobar f490( dummy[490], vec_63_bits[31], vec_63_bits[ 8] );
    foobar f491( dummy[491], vec_63_bits[32], vec_63_bits[ 8] );
    foobar f492( dummy[492], vec_63_bits[33], vec_63_bits[ 8] );
    foobar f493( dummy[493], vec_63_bits[34], vec_63_bits[ 8] );
    foobar f494( dummy[494], vec_63_bits[35], vec_63_bits[ 8] );
    foobar f495( dummy[495], vec_63_bits[36], vec_63_bits[ 8] );
    foobar f496( dummy[496], vec_63_bits[37], vec_63_bits[ 8] );
    foobar f497( dummy[497], vec_63_bits[38], vec_63_bits[ 8] );
    foobar f498( dummy[498], vec_63_bits[39], vec_63_bits[ 8] );
    foobar f499( dummy[499], vec_63_bits[40], vec_63_bits[ 8] );
    foobar f500( dummy[500], vec_63_bits[41], vec_63_bits[ 8] );
    foobar f501( dummy[501], vec_63_bits[42], vec_63_bits[ 8] );
    foobar f502( dummy[502], vec_63_bits[43], vec_63_bits[ 8] );
    foobar f503( dummy[503], vec_63_bits[44], vec_63_bits[ 8] );
    foobar f504( dummy[504], vec_63_bits[45], vec_63_bits[ 8] );
    foobar f505( dummy[505], vec_63_bits[46], vec_63_bits[ 8] );
    foobar f506( dummy[506], vec_63_bits[47], vec_63_bits[ 8] );
    foobar f507( dummy[507], vec_63_bits[48], vec_63_bits[ 8] );
    foobar f508( dummy[508], vec_63_bits[49], vec_63_bits[ 8] );
    foobar f509( dummy[509], vec_63_bits[50], vec_63_bits[ 8] );
    foobar f510( dummy[510], vec_63_bits[51], vec_63_bits[ 8] );
    foobar f511( dummy[511], vec_63_bits[52], vec_63_bits[ 8] );
    foobar f512( dummy[512], vec_63_bits[53], vec_63_bits[ 8] );
    foobar f513( dummy[513], vec_63_bits[54], vec_63_bits[ 8] );
    foobar f514( dummy[514], vec_63_bits[55], vec_63_bits[ 8] );
    foobar f515( dummy[515], vec_63_bits[56], vec_63_bits[ 8] );
    foobar f516( dummy[516], vec_63_bits[57], vec_63_bits[ 8] );
    foobar f517( dummy[517], vec_63_bits[58], vec_63_bits[ 8] );
    foobar f518( dummy[518], vec_63_bits[59], vec_63_bits[ 8] );
    foobar f519( dummy[519], vec_63_bits[60], vec_63_bits[ 8] );
    foobar f520( dummy[520], vec_63_bits[61], vec_63_bits[ 8] );
    foobar f521( dummy[521], vec_63_bits[62], vec_63_bits[ 8] );
    AN64   an8( o[8], {dummy[468], dummy[469], dummy[470], dummy[471], dummy[472], dummy[473], dummy[474], dummy[475], dummy[476], dummy[477], dummy[478], dummy[479], dummy[480], dummy[481], dummy[482], dummy[483], dummy[484], dummy[485], dummy[486], dummy[487], dummy[488], dummy[489], dummy[490], dummy[491], dummy[492], dummy[493], dummy[494], dummy[495], dummy[496], dummy[497], dummy[498], dummy[499], dummy[500], dummy[501], dummy[502], dummy[503], dummy[504], dummy[505], dummy[506], dummy[507], dummy[508], dummy[509], dummy[510], dummy[511], dummy[512], dummy[513], dummy[514], dummy[515], dummy[516], dummy[517], dummy[518], dummy[519], dummy[520], dummy[521], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f522( dummy[522], vec_63_bits[10], vec_63_bits[ 9] );
    foobar f523( dummy[523], vec_63_bits[11], vec_63_bits[ 9] );
    foobar f524( dummy[524], vec_63_bits[12], vec_63_bits[ 9] );
    foobar f525( dummy[525], vec_63_bits[13], vec_63_bits[ 9] );
    foobar f526( dummy[526], vec_63_bits[14], vec_63_bits[ 9] );
    foobar f527( dummy[527], vec_63_bits[15], vec_63_bits[ 9] );
    foobar f528( dummy[528], vec_63_bits[16], vec_63_bits[ 9] );
    foobar f529( dummy[529], vec_63_bits[17], vec_63_bits[ 9] );
    foobar f530( dummy[530], vec_63_bits[18], vec_63_bits[ 9] );
    foobar f531( dummy[531], vec_63_bits[19], vec_63_bits[ 9] );
    foobar f532( dummy[532], vec_63_bits[20], vec_63_bits[ 9] );
    foobar f533( dummy[533], vec_63_bits[21], vec_63_bits[ 9] );
    foobar f534( dummy[534], vec_63_bits[22], vec_63_bits[ 9] );
    foobar f535( dummy[535], vec_63_bits[23], vec_63_bits[ 9] );
    foobar f536( dummy[536], vec_63_bits[24], vec_63_bits[ 9] );
    foobar f537( dummy[537], vec_63_bits[25], vec_63_bits[ 9] );
    foobar f538( dummy[538], vec_63_bits[26], vec_63_bits[ 9] );
    foobar f539( dummy[539], vec_63_bits[27], vec_63_bits[ 9] );
    foobar f540( dummy[540], vec_63_bits[28], vec_63_bits[ 9] );
    foobar f541( dummy[541], vec_63_bits[29], vec_63_bits[ 9] );
    foobar f542( dummy[542], vec_63_bits[30], vec_63_bits[ 9] );
    foobar f543( dummy[543], vec_63_bits[31], vec_63_bits[ 9] );
    foobar f544( dummy[544], vec_63_bits[32], vec_63_bits[ 9] );
    foobar f545( dummy[545], vec_63_bits[33], vec_63_bits[ 9] );
    foobar f546( dummy[546], vec_63_bits[34], vec_63_bits[ 9] );
    foobar f547( dummy[547], vec_63_bits[35], vec_63_bits[ 9] );
    foobar f548( dummy[548], vec_63_bits[36], vec_63_bits[ 9] );
    foobar f549( dummy[549], vec_63_bits[37], vec_63_bits[ 9] );
    foobar f550( dummy[550], vec_63_bits[38], vec_63_bits[ 9] );
    foobar f551( dummy[551], vec_63_bits[39], vec_63_bits[ 9] );
    foobar f552( dummy[552], vec_63_bits[40], vec_63_bits[ 9] );
    foobar f553( dummy[553], vec_63_bits[41], vec_63_bits[ 9] );
    foobar f554( dummy[554], vec_63_bits[42], vec_63_bits[ 9] );
    foobar f555( dummy[555], vec_63_bits[43], vec_63_bits[ 9] );
    foobar f556( dummy[556], vec_63_bits[44], vec_63_bits[ 9] );
    foobar f557( dummy[557], vec_63_bits[45], vec_63_bits[ 9] );
    foobar f558( dummy[558], vec_63_bits[46], vec_63_bits[ 9] );
    foobar f559( dummy[559], vec_63_bits[47], vec_63_bits[ 9] );
    foobar f560( dummy[560], vec_63_bits[48], vec_63_bits[ 9] );
    foobar f561( dummy[561], vec_63_bits[49], vec_63_bits[ 9] );
    foobar f562( dummy[562], vec_63_bits[50], vec_63_bits[ 9] );
    foobar f563( dummy[563], vec_63_bits[51], vec_63_bits[ 9] );
    foobar f564( dummy[564], vec_63_bits[52], vec_63_bits[ 9] );
    foobar f565( dummy[565], vec_63_bits[53], vec_63_bits[ 9] );
    foobar f566( dummy[566], vec_63_bits[54], vec_63_bits[ 9] );
    foobar f567( dummy[567], vec_63_bits[55], vec_63_bits[ 9] );
    foobar f568( dummy[568], vec_63_bits[56], vec_63_bits[ 9] );
    foobar f569( dummy[569], vec_63_bits[57], vec_63_bits[ 9] );
    foobar f570( dummy[570], vec_63_bits[58], vec_63_bits[ 9] );
    foobar f571( dummy[571], vec_63_bits[59], vec_63_bits[ 9] );
    foobar f572( dummy[572], vec_63_bits[60], vec_63_bits[ 9] );
    foobar f573( dummy[573], vec_63_bits[61], vec_63_bits[ 9] );
    foobar f574( dummy[574], vec_63_bits[62], vec_63_bits[ 9] );
    AN64   an9( o[9], {dummy[522], dummy[523], dummy[524], dummy[525], dummy[526], dummy[527], dummy[528], dummy[529], dummy[530], dummy[531], dummy[532], dummy[533], dummy[534], dummy[535], dummy[536], dummy[537], dummy[538], dummy[539], dummy[540], dummy[541], dummy[542], dummy[543], dummy[544], dummy[545], dummy[546], dummy[547], dummy[548], dummy[549], dummy[550], dummy[551], dummy[552], dummy[553], dummy[554], dummy[555], dummy[556], dummy[557], dummy[558], dummy[559], dummy[560], dummy[561], dummy[562], dummy[563], dummy[564], dummy[565], dummy[566], dummy[567], dummy[568], dummy[569], dummy[570], dummy[571], dummy[572], dummy[573], dummy[574], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f575( dummy[575], vec_63_bits[11], vec_63_bits[10] );
    foobar f576( dummy[576], vec_63_bits[12], vec_63_bits[10] );
    foobar f577( dummy[577], vec_63_bits[13], vec_63_bits[10] );
    foobar f578( dummy[578], vec_63_bits[14], vec_63_bits[10] );
    foobar f579( dummy[579], vec_63_bits[15], vec_63_bits[10] );
    foobar f580( dummy[580], vec_63_bits[16], vec_63_bits[10] );
    foobar f581( dummy[581], vec_63_bits[17], vec_63_bits[10] );
    foobar f582( dummy[582], vec_63_bits[18], vec_63_bits[10] );
    foobar f583( dummy[583], vec_63_bits[19], vec_63_bits[10] );
    foobar f584( dummy[584], vec_63_bits[20], vec_63_bits[10] );
    foobar f585( dummy[585], vec_63_bits[21], vec_63_bits[10] );
    foobar f586( dummy[586], vec_63_bits[22], vec_63_bits[10] );
    foobar f587( dummy[587], vec_63_bits[23], vec_63_bits[10] );
    foobar f588( dummy[588], vec_63_bits[24], vec_63_bits[10] );
    foobar f589( dummy[589], vec_63_bits[25], vec_63_bits[10] );
    foobar f590( dummy[590], vec_63_bits[26], vec_63_bits[10] );
    foobar f591( dummy[591], vec_63_bits[27], vec_63_bits[10] );
    foobar f592( dummy[592], vec_63_bits[28], vec_63_bits[10] );
    foobar f593( dummy[593], vec_63_bits[29], vec_63_bits[10] );
    foobar f594( dummy[594], vec_63_bits[30], vec_63_bits[10] );
    foobar f595( dummy[595], vec_63_bits[31], vec_63_bits[10] );
    foobar f596( dummy[596], vec_63_bits[32], vec_63_bits[10] );
    foobar f597( dummy[597], vec_63_bits[33], vec_63_bits[10] );
    foobar f598( dummy[598], vec_63_bits[34], vec_63_bits[10] );
    foobar f599( dummy[599], vec_63_bits[35], vec_63_bits[10] );
    foobar f600( dummy[600], vec_63_bits[36], vec_63_bits[10] );
    foobar f601( dummy[601], vec_63_bits[37], vec_63_bits[10] );
    foobar f602( dummy[602], vec_63_bits[38], vec_63_bits[10] );
    foobar f603( dummy[603], vec_63_bits[39], vec_63_bits[10] );
    foobar f604( dummy[604], vec_63_bits[40], vec_63_bits[10] );
    foobar f605( dummy[605], vec_63_bits[41], vec_63_bits[10] );
    foobar f606( dummy[606], vec_63_bits[42], vec_63_bits[10] );
    foobar f607( dummy[607], vec_63_bits[43], vec_63_bits[10] );
    foobar f608( dummy[608], vec_63_bits[44], vec_63_bits[10] );
    foobar f609( dummy[609], vec_63_bits[45], vec_63_bits[10] );
    foobar f610( dummy[610], vec_63_bits[46], vec_63_bits[10] );
    foobar f611( dummy[611], vec_63_bits[47], vec_63_bits[10] );
    foobar f612( dummy[612], vec_63_bits[48], vec_63_bits[10] );
    foobar f613( dummy[613], vec_63_bits[49], vec_63_bits[10] );
    foobar f614( dummy[614], vec_63_bits[50], vec_63_bits[10] );
    foobar f615( dummy[615], vec_63_bits[51], vec_63_bits[10] );
    foobar f616( dummy[616], vec_63_bits[52], vec_63_bits[10] );
    foobar f617( dummy[617], vec_63_bits[53], vec_63_bits[10] );
    foobar f618( dummy[618], vec_63_bits[54], vec_63_bits[10] );
    foobar f619( dummy[619], vec_63_bits[55], vec_63_bits[10] );
    foobar f620( dummy[620], vec_63_bits[56], vec_63_bits[10] );
    foobar f621( dummy[621], vec_63_bits[57], vec_63_bits[10] );
    foobar f622( dummy[622], vec_63_bits[58], vec_63_bits[10] );
    foobar f623( dummy[623], vec_63_bits[59], vec_63_bits[10] );
    foobar f624( dummy[624], vec_63_bits[60], vec_63_bits[10] );
    foobar f625( dummy[625], vec_63_bits[61], vec_63_bits[10] );
    foobar f626( dummy[626], vec_63_bits[62], vec_63_bits[10] );
    AN64   an10( o[10], {dummy[575], dummy[576], dummy[577], dummy[578], dummy[579], dummy[580], dummy[581], dummy[582], dummy[583], dummy[584], dummy[585], dummy[586], dummy[587], dummy[588], dummy[589], dummy[590], dummy[591], dummy[592], dummy[593], dummy[594], dummy[595], dummy[596], dummy[597], dummy[598], dummy[599], dummy[600], dummy[601], dummy[602], dummy[603], dummy[604], dummy[605], dummy[606], dummy[607], dummy[608], dummy[609], dummy[610], dummy[611], dummy[612], dummy[613], dummy[614], dummy[615], dummy[616], dummy[617], dummy[618], dummy[619], dummy[620], dummy[621], dummy[622], dummy[623], dummy[624], dummy[625], dummy[626], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f627( dummy[627], vec_63_bits[12], vec_63_bits[11] );
    foobar f628( dummy[628], vec_63_bits[13], vec_63_bits[11] );
    foobar f629( dummy[629], vec_63_bits[14], vec_63_bits[11] );
    foobar f630( dummy[630], vec_63_bits[15], vec_63_bits[11] );
    foobar f631( dummy[631], vec_63_bits[16], vec_63_bits[11] );
    foobar f632( dummy[632], vec_63_bits[17], vec_63_bits[11] );
    foobar f633( dummy[633], vec_63_bits[18], vec_63_bits[11] );
    foobar f634( dummy[634], vec_63_bits[19], vec_63_bits[11] );
    foobar f635( dummy[635], vec_63_bits[20], vec_63_bits[11] );
    foobar f636( dummy[636], vec_63_bits[21], vec_63_bits[11] );
    foobar f637( dummy[637], vec_63_bits[22], vec_63_bits[11] );
    foobar f638( dummy[638], vec_63_bits[23], vec_63_bits[11] );
    foobar f639( dummy[639], vec_63_bits[24], vec_63_bits[11] );
    foobar f640( dummy[640], vec_63_bits[25], vec_63_bits[11] );
    foobar f641( dummy[641], vec_63_bits[26], vec_63_bits[11] );
    foobar f642( dummy[642], vec_63_bits[27], vec_63_bits[11] );
    foobar f643( dummy[643], vec_63_bits[28], vec_63_bits[11] );
    foobar f644( dummy[644], vec_63_bits[29], vec_63_bits[11] );
    foobar f645( dummy[645], vec_63_bits[30], vec_63_bits[11] );
    foobar f646( dummy[646], vec_63_bits[31], vec_63_bits[11] );
    foobar f647( dummy[647], vec_63_bits[32], vec_63_bits[11] );
    foobar f648( dummy[648], vec_63_bits[33], vec_63_bits[11] );
    foobar f649( dummy[649], vec_63_bits[34], vec_63_bits[11] );
    foobar f650( dummy[650], vec_63_bits[35], vec_63_bits[11] );
    foobar f651( dummy[651], vec_63_bits[36], vec_63_bits[11] );
    foobar f652( dummy[652], vec_63_bits[37], vec_63_bits[11] );
    foobar f653( dummy[653], vec_63_bits[38], vec_63_bits[11] );
    foobar f654( dummy[654], vec_63_bits[39], vec_63_bits[11] );
    foobar f655( dummy[655], vec_63_bits[40], vec_63_bits[11] );
    foobar f656( dummy[656], vec_63_bits[41], vec_63_bits[11] );
    foobar f657( dummy[657], vec_63_bits[42], vec_63_bits[11] );
    foobar f658( dummy[658], vec_63_bits[43], vec_63_bits[11] );
    foobar f659( dummy[659], vec_63_bits[44], vec_63_bits[11] );
    foobar f660( dummy[660], vec_63_bits[45], vec_63_bits[11] );
    foobar f661( dummy[661], vec_63_bits[46], vec_63_bits[11] );
    foobar f662( dummy[662], vec_63_bits[47], vec_63_bits[11] );
    foobar f663( dummy[663], vec_63_bits[48], vec_63_bits[11] );
    foobar f664( dummy[664], vec_63_bits[49], vec_63_bits[11] );
    foobar f665( dummy[665], vec_63_bits[50], vec_63_bits[11] );
    foobar f666( dummy[666], vec_63_bits[51], vec_63_bits[11] );
    foobar f667( dummy[667], vec_63_bits[52], vec_63_bits[11] );
    foobar f668( dummy[668], vec_63_bits[53], vec_63_bits[11] );
    foobar f669( dummy[669], vec_63_bits[54], vec_63_bits[11] );
    foobar f670( dummy[670], vec_63_bits[55], vec_63_bits[11] );
    foobar f671( dummy[671], vec_63_bits[56], vec_63_bits[11] );
    foobar f672( dummy[672], vec_63_bits[57], vec_63_bits[11] );
    foobar f673( dummy[673], vec_63_bits[58], vec_63_bits[11] );
    foobar f674( dummy[674], vec_63_bits[59], vec_63_bits[11] );
    foobar f675( dummy[675], vec_63_bits[60], vec_63_bits[11] );
    foobar f676( dummy[676], vec_63_bits[61], vec_63_bits[11] );
    foobar f677( dummy[677], vec_63_bits[62], vec_63_bits[11] );
    AN64   an11( o[11], {dummy[627], dummy[628], dummy[629], dummy[630], dummy[631], dummy[632], dummy[633], dummy[634], dummy[635], dummy[636], dummy[637], dummy[638], dummy[639], dummy[640], dummy[641], dummy[642], dummy[643], dummy[644], dummy[645], dummy[646], dummy[647], dummy[648], dummy[649], dummy[650], dummy[651], dummy[652], dummy[653], dummy[654], dummy[655], dummy[656], dummy[657], dummy[658], dummy[659], dummy[660], dummy[661], dummy[662], dummy[663], dummy[664], dummy[665], dummy[666], dummy[667], dummy[668], dummy[669], dummy[670], dummy[671], dummy[672], dummy[673], dummy[674], dummy[675], dummy[676], dummy[677], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f678( dummy[678], vec_63_bits[13], vec_63_bits[12] );
    foobar f679( dummy[679], vec_63_bits[14], vec_63_bits[12] );
    foobar f680( dummy[680], vec_63_bits[15], vec_63_bits[12] );
    foobar f681( dummy[681], vec_63_bits[16], vec_63_bits[12] );
    foobar f682( dummy[682], vec_63_bits[17], vec_63_bits[12] );
    foobar f683( dummy[683], vec_63_bits[18], vec_63_bits[12] );
    foobar f684( dummy[684], vec_63_bits[19], vec_63_bits[12] );
    foobar f685( dummy[685], vec_63_bits[20], vec_63_bits[12] );
    foobar f686( dummy[686], vec_63_bits[21], vec_63_bits[12] );
    foobar f687( dummy[687], vec_63_bits[22], vec_63_bits[12] );
    foobar f688( dummy[688], vec_63_bits[23], vec_63_bits[12] );
    foobar f689( dummy[689], vec_63_bits[24], vec_63_bits[12] );
    foobar f690( dummy[690], vec_63_bits[25], vec_63_bits[12] );
    foobar f691( dummy[691], vec_63_bits[26], vec_63_bits[12] );
    foobar f692( dummy[692], vec_63_bits[27], vec_63_bits[12] );
    foobar f693( dummy[693], vec_63_bits[28], vec_63_bits[12] );
    foobar f694( dummy[694], vec_63_bits[29], vec_63_bits[12] );
    foobar f695( dummy[695], vec_63_bits[30], vec_63_bits[12] );
    foobar f696( dummy[696], vec_63_bits[31], vec_63_bits[12] );
    foobar f697( dummy[697], vec_63_bits[32], vec_63_bits[12] );
    foobar f698( dummy[698], vec_63_bits[33], vec_63_bits[12] );
    foobar f699( dummy[699], vec_63_bits[34], vec_63_bits[12] );
    foobar f700( dummy[700], vec_63_bits[35], vec_63_bits[12] );
    foobar f701( dummy[701], vec_63_bits[36], vec_63_bits[12] );
    foobar f702( dummy[702], vec_63_bits[37], vec_63_bits[12] );
    foobar f703( dummy[703], vec_63_bits[38], vec_63_bits[12] );
    foobar f704( dummy[704], vec_63_bits[39], vec_63_bits[12] );
    foobar f705( dummy[705], vec_63_bits[40], vec_63_bits[12] );
    foobar f706( dummy[706], vec_63_bits[41], vec_63_bits[12] );
    foobar f707( dummy[707], vec_63_bits[42], vec_63_bits[12] );
    foobar f708( dummy[708], vec_63_bits[43], vec_63_bits[12] );
    foobar f709( dummy[709], vec_63_bits[44], vec_63_bits[12] );
    foobar f710( dummy[710], vec_63_bits[45], vec_63_bits[12] );
    foobar f711( dummy[711], vec_63_bits[46], vec_63_bits[12] );
    foobar f712( dummy[712], vec_63_bits[47], vec_63_bits[12] );
    foobar f713( dummy[713], vec_63_bits[48], vec_63_bits[12] );
    foobar f714( dummy[714], vec_63_bits[49], vec_63_bits[12] );
    foobar f715( dummy[715], vec_63_bits[50], vec_63_bits[12] );
    foobar f716( dummy[716], vec_63_bits[51], vec_63_bits[12] );
    foobar f717( dummy[717], vec_63_bits[52], vec_63_bits[12] );
    foobar f718( dummy[718], vec_63_bits[53], vec_63_bits[12] );
    foobar f719( dummy[719], vec_63_bits[54], vec_63_bits[12] );
    foobar f720( dummy[720], vec_63_bits[55], vec_63_bits[12] );
    foobar f721( dummy[721], vec_63_bits[56], vec_63_bits[12] );
    foobar f722( dummy[722], vec_63_bits[57], vec_63_bits[12] );
    foobar f723( dummy[723], vec_63_bits[58], vec_63_bits[12] );
    foobar f724( dummy[724], vec_63_bits[59], vec_63_bits[12] );
    foobar f725( dummy[725], vec_63_bits[60], vec_63_bits[12] );
    foobar f726( dummy[726], vec_63_bits[61], vec_63_bits[12] );
    foobar f727( dummy[727], vec_63_bits[62], vec_63_bits[12] );
    AN64   an12( o[12], {dummy[678], dummy[679], dummy[680], dummy[681], dummy[682], dummy[683], dummy[684], dummy[685], dummy[686], dummy[687], dummy[688], dummy[689], dummy[690], dummy[691], dummy[692], dummy[693], dummy[694], dummy[695], dummy[696], dummy[697], dummy[698], dummy[699], dummy[700], dummy[701], dummy[702], dummy[703], dummy[704], dummy[705], dummy[706], dummy[707], dummy[708], dummy[709], dummy[710], dummy[711], dummy[712], dummy[713], dummy[714], dummy[715], dummy[716], dummy[717], dummy[718], dummy[719], dummy[720], dummy[721], dummy[722], dummy[723], dummy[724], dummy[725], dummy[726], dummy[727], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f728( dummy[728], vec_63_bits[14], vec_63_bits[13] );
    foobar f729( dummy[729], vec_63_bits[15], vec_63_bits[13] );
    foobar f730( dummy[730], vec_63_bits[16], vec_63_bits[13] );
    foobar f731( dummy[731], vec_63_bits[17], vec_63_bits[13] );
    foobar f732( dummy[732], vec_63_bits[18], vec_63_bits[13] );
    foobar f733( dummy[733], vec_63_bits[19], vec_63_bits[13] );
    foobar f734( dummy[734], vec_63_bits[20], vec_63_bits[13] );
    foobar f735( dummy[735], vec_63_bits[21], vec_63_bits[13] );
    foobar f736( dummy[736], vec_63_bits[22], vec_63_bits[13] );
    foobar f737( dummy[737], vec_63_bits[23], vec_63_bits[13] );
    foobar f738( dummy[738], vec_63_bits[24], vec_63_bits[13] );
    foobar f739( dummy[739], vec_63_bits[25], vec_63_bits[13] );
    foobar f740( dummy[740], vec_63_bits[26], vec_63_bits[13] );
    foobar f741( dummy[741], vec_63_bits[27], vec_63_bits[13] );
    foobar f742( dummy[742], vec_63_bits[28], vec_63_bits[13] );
    foobar f743( dummy[743], vec_63_bits[29], vec_63_bits[13] );
    foobar f744( dummy[744], vec_63_bits[30], vec_63_bits[13] );
    foobar f745( dummy[745], vec_63_bits[31], vec_63_bits[13] );
    foobar f746( dummy[746], vec_63_bits[32], vec_63_bits[13] );
    foobar f747( dummy[747], vec_63_bits[33], vec_63_bits[13] );
    foobar f748( dummy[748], vec_63_bits[34], vec_63_bits[13] );
    foobar f749( dummy[749], vec_63_bits[35], vec_63_bits[13] );
    foobar f750( dummy[750], vec_63_bits[36], vec_63_bits[13] );
    foobar f751( dummy[751], vec_63_bits[37], vec_63_bits[13] );
    foobar f752( dummy[752], vec_63_bits[38], vec_63_bits[13] );
    foobar f753( dummy[753], vec_63_bits[39], vec_63_bits[13] );
    foobar f754( dummy[754], vec_63_bits[40], vec_63_bits[13] );
    foobar f755( dummy[755], vec_63_bits[41], vec_63_bits[13] );
    foobar f756( dummy[756], vec_63_bits[42], vec_63_bits[13] );
    foobar f757( dummy[757], vec_63_bits[43], vec_63_bits[13] );
    foobar f758( dummy[758], vec_63_bits[44], vec_63_bits[13] );
    foobar f759( dummy[759], vec_63_bits[45], vec_63_bits[13] );
    foobar f760( dummy[760], vec_63_bits[46], vec_63_bits[13] );
    foobar f761( dummy[761], vec_63_bits[47], vec_63_bits[13] );
    foobar f762( dummy[762], vec_63_bits[48], vec_63_bits[13] );
    foobar f763( dummy[763], vec_63_bits[49], vec_63_bits[13] );
    foobar f764( dummy[764], vec_63_bits[50], vec_63_bits[13] );
    foobar f765( dummy[765], vec_63_bits[51], vec_63_bits[13] );
    foobar f766( dummy[766], vec_63_bits[52], vec_63_bits[13] );
    foobar f767( dummy[767], vec_63_bits[53], vec_63_bits[13] );
    foobar f768( dummy[768], vec_63_bits[54], vec_63_bits[13] );
    foobar f769( dummy[769], vec_63_bits[55], vec_63_bits[13] );
    foobar f770( dummy[770], vec_63_bits[56], vec_63_bits[13] );
    foobar f771( dummy[771], vec_63_bits[57], vec_63_bits[13] );
    foobar f772( dummy[772], vec_63_bits[58], vec_63_bits[13] );
    foobar f773( dummy[773], vec_63_bits[59], vec_63_bits[13] );
    foobar f774( dummy[774], vec_63_bits[60], vec_63_bits[13] );
    foobar f775( dummy[775], vec_63_bits[61], vec_63_bits[13] );
    foobar f776( dummy[776], vec_63_bits[62], vec_63_bits[13] );
    AN64   an13( o[13], {dummy[728], dummy[729], dummy[730], dummy[731], dummy[732], dummy[733], dummy[734], dummy[735], dummy[736], dummy[737], dummy[738], dummy[739], dummy[740], dummy[741], dummy[742], dummy[743], dummy[744], dummy[745], dummy[746], dummy[747], dummy[748], dummy[749], dummy[750], dummy[751], dummy[752], dummy[753], dummy[754], dummy[755], dummy[756], dummy[757], dummy[758], dummy[759], dummy[760], dummy[761], dummy[762], dummy[763], dummy[764], dummy[765], dummy[766], dummy[767], dummy[768], dummy[769], dummy[770], dummy[771], dummy[772], dummy[773], dummy[774], dummy[775], dummy[776], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f777( dummy[777], vec_63_bits[15], vec_63_bits[14] );
    foobar f778( dummy[778], vec_63_bits[16], vec_63_bits[14] );
    foobar f779( dummy[779], vec_63_bits[17], vec_63_bits[14] );
    foobar f780( dummy[780], vec_63_bits[18], vec_63_bits[14] );
    foobar f781( dummy[781], vec_63_bits[19], vec_63_bits[14] );
    foobar f782( dummy[782], vec_63_bits[20], vec_63_bits[14] );
    foobar f783( dummy[783], vec_63_bits[21], vec_63_bits[14] );
    foobar f784( dummy[784], vec_63_bits[22], vec_63_bits[14] );
    foobar f785( dummy[785], vec_63_bits[23], vec_63_bits[14] );
    foobar f786( dummy[786], vec_63_bits[24], vec_63_bits[14] );
    foobar f787( dummy[787], vec_63_bits[25], vec_63_bits[14] );
    foobar f788( dummy[788], vec_63_bits[26], vec_63_bits[14] );
    foobar f789( dummy[789], vec_63_bits[27], vec_63_bits[14] );
    foobar f790( dummy[790], vec_63_bits[28], vec_63_bits[14] );
    foobar f791( dummy[791], vec_63_bits[29], vec_63_bits[14] );
    foobar f792( dummy[792], vec_63_bits[30], vec_63_bits[14] );
    foobar f793( dummy[793], vec_63_bits[31], vec_63_bits[14] );
    foobar f794( dummy[794], vec_63_bits[32], vec_63_bits[14] );
    foobar f795( dummy[795], vec_63_bits[33], vec_63_bits[14] );
    foobar f796( dummy[796], vec_63_bits[34], vec_63_bits[14] );
    foobar f797( dummy[797], vec_63_bits[35], vec_63_bits[14] );
    foobar f798( dummy[798], vec_63_bits[36], vec_63_bits[14] );
    foobar f799( dummy[799], vec_63_bits[37], vec_63_bits[14] );
    foobar f800( dummy[800], vec_63_bits[38], vec_63_bits[14] );
    foobar f801( dummy[801], vec_63_bits[39], vec_63_bits[14] );
    foobar f802( dummy[802], vec_63_bits[40], vec_63_bits[14] );
    foobar f803( dummy[803], vec_63_bits[41], vec_63_bits[14] );
    foobar f804( dummy[804], vec_63_bits[42], vec_63_bits[14] );
    foobar f805( dummy[805], vec_63_bits[43], vec_63_bits[14] );
    foobar f806( dummy[806], vec_63_bits[44], vec_63_bits[14] );
    foobar f807( dummy[807], vec_63_bits[45], vec_63_bits[14] );
    foobar f808( dummy[808], vec_63_bits[46], vec_63_bits[14] );
    foobar f809( dummy[809], vec_63_bits[47], vec_63_bits[14] );
    foobar f810( dummy[810], vec_63_bits[48], vec_63_bits[14] );
    foobar f811( dummy[811], vec_63_bits[49], vec_63_bits[14] );
    foobar f812( dummy[812], vec_63_bits[50], vec_63_bits[14] );
    foobar f813( dummy[813], vec_63_bits[51], vec_63_bits[14] );
    foobar f814( dummy[814], vec_63_bits[52], vec_63_bits[14] );
    foobar f815( dummy[815], vec_63_bits[53], vec_63_bits[14] );
    foobar f816( dummy[816], vec_63_bits[54], vec_63_bits[14] );
    foobar f817( dummy[817], vec_63_bits[55], vec_63_bits[14] );
    foobar f818( dummy[818], vec_63_bits[56], vec_63_bits[14] );
    foobar f819( dummy[819], vec_63_bits[57], vec_63_bits[14] );
    foobar f820( dummy[820], vec_63_bits[58], vec_63_bits[14] );
    foobar f821( dummy[821], vec_63_bits[59], vec_63_bits[14] );
    foobar f822( dummy[822], vec_63_bits[60], vec_63_bits[14] );
    foobar f823( dummy[823], vec_63_bits[61], vec_63_bits[14] );
    foobar f824( dummy[824], vec_63_bits[62], vec_63_bits[14] );
    AN64   an14( o[14], {dummy[777], dummy[778], dummy[779], dummy[780], dummy[781], dummy[782], dummy[783], dummy[784], dummy[785], dummy[786], dummy[787], dummy[788], dummy[789], dummy[790], dummy[791], dummy[792], dummy[793], dummy[794], dummy[795], dummy[796], dummy[797], dummy[798], dummy[799], dummy[800], dummy[801], dummy[802], dummy[803], dummy[804], dummy[805], dummy[806], dummy[807], dummy[808], dummy[809], dummy[810], dummy[811], dummy[812], dummy[813], dummy[814], dummy[815], dummy[816], dummy[817], dummy[818], dummy[819], dummy[820], dummy[821], dummy[822], dummy[823], dummy[824], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f825( dummy[825], vec_63_bits[16], vec_63_bits[15] );
    foobar f826( dummy[826], vec_63_bits[17], vec_63_bits[15] );
    foobar f827( dummy[827], vec_63_bits[18], vec_63_bits[15] );
    foobar f828( dummy[828], vec_63_bits[19], vec_63_bits[15] );
    foobar f829( dummy[829], vec_63_bits[20], vec_63_bits[15] );
    foobar f830( dummy[830], vec_63_bits[21], vec_63_bits[15] );
    foobar f831( dummy[831], vec_63_bits[22], vec_63_bits[15] );
    foobar f832( dummy[832], vec_63_bits[23], vec_63_bits[15] );
    foobar f833( dummy[833], vec_63_bits[24], vec_63_bits[15] );
    foobar f834( dummy[834], vec_63_bits[25], vec_63_bits[15] );
    foobar f835( dummy[835], vec_63_bits[26], vec_63_bits[15] );
    foobar f836( dummy[836], vec_63_bits[27], vec_63_bits[15] );
    foobar f837( dummy[837], vec_63_bits[28], vec_63_bits[15] );
    foobar f838( dummy[838], vec_63_bits[29], vec_63_bits[15] );
    foobar f839( dummy[839], vec_63_bits[30], vec_63_bits[15] );
    foobar f840( dummy[840], vec_63_bits[31], vec_63_bits[15] );
    foobar f841( dummy[841], vec_63_bits[32], vec_63_bits[15] );
    foobar f842( dummy[842], vec_63_bits[33], vec_63_bits[15] );
    foobar f843( dummy[843], vec_63_bits[34], vec_63_bits[15] );
    foobar f844( dummy[844], vec_63_bits[35], vec_63_bits[15] );
    foobar f845( dummy[845], vec_63_bits[36], vec_63_bits[15] );
    foobar f846( dummy[846], vec_63_bits[37], vec_63_bits[15] );
    foobar f847( dummy[847], vec_63_bits[38], vec_63_bits[15] );
    foobar f848( dummy[848], vec_63_bits[39], vec_63_bits[15] );
    foobar f849( dummy[849], vec_63_bits[40], vec_63_bits[15] );
    foobar f850( dummy[850], vec_63_bits[41], vec_63_bits[15] );
    foobar f851( dummy[851], vec_63_bits[42], vec_63_bits[15] );
    foobar f852( dummy[852], vec_63_bits[43], vec_63_bits[15] );
    foobar f853( dummy[853], vec_63_bits[44], vec_63_bits[15] );
    foobar f854( dummy[854], vec_63_bits[45], vec_63_bits[15] );
    foobar f855( dummy[855], vec_63_bits[46], vec_63_bits[15] );
    foobar f856( dummy[856], vec_63_bits[47], vec_63_bits[15] );
    foobar f857( dummy[857], vec_63_bits[48], vec_63_bits[15] );
    foobar f858( dummy[858], vec_63_bits[49], vec_63_bits[15] );
    foobar f859( dummy[859], vec_63_bits[50], vec_63_bits[15] );
    foobar f860( dummy[860], vec_63_bits[51], vec_63_bits[15] );
    foobar f861( dummy[861], vec_63_bits[52], vec_63_bits[15] );
    foobar f862( dummy[862], vec_63_bits[53], vec_63_bits[15] );
    foobar f863( dummy[863], vec_63_bits[54], vec_63_bits[15] );
    foobar f864( dummy[864], vec_63_bits[55], vec_63_bits[15] );
    foobar f865( dummy[865], vec_63_bits[56], vec_63_bits[15] );
    foobar f866( dummy[866], vec_63_bits[57], vec_63_bits[15] );
    foobar f867( dummy[867], vec_63_bits[58], vec_63_bits[15] );
    foobar f868( dummy[868], vec_63_bits[59], vec_63_bits[15] );
    foobar f869( dummy[869], vec_63_bits[60], vec_63_bits[15] );
    foobar f870( dummy[870], vec_63_bits[61], vec_63_bits[15] );
    foobar f871( dummy[871], vec_63_bits[62], vec_63_bits[15] );
    AN64   an15( o[15], {dummy[825], dummy[826], dummy[827], dummy[828], dummy[829], dummy[830], dummy[831], dummy[832], dummy[833], dummy[834], dummy[835], dummy[836], dummy[837], dummy[838], dummy[839], dummy[840], dummy[841], dummy[842], dummy[843], dummy[844], dummy[845], dummy[846], dummy[847], dummy[848], dummy[849], dummy[850], dummy[851], dummy[852], dummy[853], dummy[854], dummy[855], dummy[856], dummy[857], dummy[858], dummy[859], dummy[860], dummy[861], dummy[862], dummy[863], dummy[864], dummy[865], dummy[866], dummy[867], dummy[868], dummy[869], dummy[870], dummy[871], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f872( dummy[872], vec_63_bits[17], vec_63_bits[16] );
    foobar f873( dummy[873], vec_63_bits[18], vec_63_bits[16] );
    foobar f874( dummy[874], vec_63_bits[19], vec_63_bits[16] );
    foobar f875( dummy[875], vec_63_bits[20], vec_63_bits[16] );
    foobar f876( dummy[876], vec_63_bits[21], vec_63_bits[16] );
    foobar f877( dummy[877], vec_63_bits[22], vec_63_bits[16] );
    foobar f878( dummy[878], vec_63_bits[23], vec_63_bits[16] );
    foobar f879( dummy[879], vec_63_bits[24], vec_63_bits[16] );
    foobar f880( dummy[880], vec_63_bits[25], vec_63_bits[16] );
    foobar f881( dummy[881], vec_63_bits[26], vec_63_bits[16] );
    foobar f882( dummy[882], vec_63_bits[27], vec_63_bits[16] );
    foobar f883( dummy[883], vec_63_bits[28], vec_63_bits[16] );
    foobar f884( dummy[884], vec_63_bits[29], vec_63_bits[16] );
    foobar f885( dummy[885], vec_63_bits[30], vec_63_bits[16] );
    foobar f886( dummy[886], vec_63_bits[31], vec_63_bits[16] );
    foobar f887( dummy[887], vec_63_bits[32], vec_63_bits[16] );
    foobar f888( dummy[888], vec_63_bits[33], vec_63_bits[16] );
    foobar f889( dummy[889], vec_63_bits[34], vec_63_bits[16] );
    foobar f890( dummy[890], vec_63_bits[35], vec_63_bits[16] );
    foobar f891( dummy[891], vec_63_bits[36], vec_63_bits[16] );
    foobar f892( dummy[892], vec_63_bits[37], vec_63_bits[16] );
    foobar f893( dummy[893], vec_63_bits[38], vec_63_bits[16] );
    foobar f894( dummy[894], vec_63_bits[39], vec_63_bits[16] );
    foobar f895( dummy[895], vec_63_bits[40], vec_63_bits[16] );
    foobar f896( dummy[896], vec_63_bits[41], vec_63_bits[16] );
    foobar f897( dummy[897], vec_63_bits[42], vec_63_bits[16] );
    foobar f898( dummy[898], vec_63_bits[43], vec_63_bits[16] );
    foobar f899( dummy[899], vec_63_bits[44], vec_63_bits[16] );
    foobar f900( dummy[900], vec_63_bits[45], vec_63_bits[16] );
    foobar f901( dummy[901], vec_63_bits[46], vec_63_bits[16] );
    foobar f902( dummy[902], vec_63_bits[47], vec_63_bits[16] );
    foobar f903( dummy[903], vec_63_bits[48], vec_63_bits[16] );
    foobar f904( dummy[904], vec_63_bits[49], vec_63_bits[16] );
    foobar f905( dummy[905], vec_63_bits[50], vec_63_bits[16] );
    foobar f906( dummy[906], vec_63_bits[51], vec_63_bits[16] );
    foobar f907( dummy[907], vec_63_bits[52], vec_63_bits[16] );
    foobar f908( dummy[908], vec_63_bits[53], vec_63_bits[16] );
    foobar f909( dummy[909], vec_63_bits[54], vec_63_bits[16] );
    foobar f910( dummy[910], vec_63_bits[55], vec_63_bits[16] );
    foobar f911( dummy[911], vec_63_bits[56], vec_63_bits[16] );
    foobar f912( dummy[912], vec_63_bits[57], vec_63_bits[16] );
    foobar f913( dummy[913], vec_63_bits[58], vec_63_bits[16] );
    foobar f914( dummy[914], vec_63_bits[59], vec_63_bits[16] );
    foobar f915( dummy[915], vec_63_bits[60], vec_63_bits[16] );
    foobar f916( dummy[916], vec_63_bits[61], vec_63_bits[16] );
    foobar f917( dummy[917], vec_63_bits[62], vec_63_bits[16] );
    AN64   an16( o[16], {dummy[872], dummy[873], dummy[874], dummy[875], dummy[876], dummy[877], dummy[878], dummy[879], dummy[880], dummy[881], dummy[882], dummy[883], dummy[884], dummy[885], dummy[886], dummy[887], dummy[888], dummy[889], dummy[890], dummy[891], dummy[892], dummy[893], dummy[894], dummy[895], dummy[896], dummy[897], dummy[898], dummy[899], dummy[900], dummy[901], dummy[902], dummy[903], dummy[904], dummy[905], dummy[906], dummy[907], dummy[908], dummy[909], dummy[910], dummy[911], dummy[912], dummy[913], dummy[914], dummy[915], dummy[916], dummy[917], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f918( dummy[918], vec_63_bits[18], vec_63_bits[17] );
    foobar f919( dummy[919], vec_63_bits[19], vec_63_bits[17] );
    foobar f920( dummy[920], vec_63_bits[20], vec_63_bits[17] );
    foobar f921( dummy[921], vec_63_bits[21], vec_63_bits[17] );
    foobar f922( dummy[922], vec_63_bits[22], vec_63_bits[17] );
    foobar f923( dummy[923], vec_63_bits[23], vec_63_bits[17] );
    foobar f924( dummy[924], vec_63_bits[24], vec_63_bits[17] );
    foobar f925( dummy[925], vec_63_bits[25], vec_63_bits[17] );
    foobar f926( dummy[926], vec_63_bits[26], vec_63_bits[17] );
    foobar f927( dummy[927], vec_63_bits[27], vec_63_bits[17] );
    foobar f928( dummy[928], vec_63_bits[28], vec_63_bits[17] );
    foobar f929( dummy[929], vec_63_bits[29], vec_63_bits[17] );
    foobar f930( dummy[930], vec_63_bits[30], vec_63_bits[17] );
    foobar f931( dummy[931], vec_63_bits[31], vec_63_bits[17] );
    foobar f932( dummy[932], vec_63_bits[32], vec_63_bits[17] );
    foobar f933( dummy[933], vec_63_bits[33], vec_63_bits[17] );
    foobar f934( dummy[934], vec_63_bits[34], vec_63_bits[17] );
    foobar f935( dummy[935], vec_63_bits[35], vec_63_bits[17] );
    foobar f936( dummy[936], vec_63_bits[36], vec_63_bits[17] );
    foobar f937( dummy[937], vec_63_bits[37], vec_63_bits[17] );
    foobar f938( dummy[938], vec_63_bits[38], vec_63_bits[17] );
    foobar f939( dummy[939], vec_63_bits[39], vec_63_bits[17] );
    foobar f940( dummy[940], vec_63_bits[40], vec_63_bits[17] );
    foobar f941( dummy[941], vec_63_bits[41], vec_63_bits[17] );
    foobar f942( dummy[942], vec_63_bits[42], vec_63_bits[17] );
    foobar f943( dummy[943], vec_63_bits[43], vec_63_bits[17] );
    foobar f944( dummy[944], vec_63_bits[44], vec_63_bits[17] );
    foobar f945( dummy[945], vec_63_bits[45], vec_63_bits[17] );
    foobar f946( dummy[946], vec_63_bits[46], vec_63_bits[17] );
    foobar f947( dummy[947], vec_63_bits[47], vec_63_bits[17] );
    foobar f948( dummy[948], vec_63_bits[48], vec_63_bits[17] );
    foobar f949( dummy[949], vec_63_bits[49], vec_63_bits[17] );
    foobar f950( dummy[950], vec_63_bits[50], vec_63_bits[17] );
    foobar f951( dummy[951], vec_63_bits[51], vec_63_bits[17] );
    foobar f952( dummy[952], vec_63_bits[52], vec_63_bits[17] );
    foobar f953( dummy[953], vec_63_bits[53], vec_63_bits[17] );
    foobar f954( dummy[954], vec_63_bits[54], vec_63_bits[17] );
    foobar f955( dummy[955], vec_63_bits[55], vec_63_bits[17] );
    foobar f956( dummy[956], vec_63_bits[56], vec_63_bits[17] );
    foobar f957( dummy[957], vec_63_bits[57], vec_63_bits[17] );
    foobar f958( dummy[958], vec_63_bits[58], vec_63_bits[17] );
    foobar f959( dummy[959], vec_63_bits[59], vec_63_bits[17] );
    foobar f960( dummy[960], vec_63_bits[60], vec_63_bits[17] );
    foobar f961( dummy[961], vec_63_bits[61], vec_63_bits[17] );
    foobar f962( dummy[962], vec_63_bits[62], vec_63_bits[17] );
    AN64   an17( o[17], {dummy[918], dummy[919], dummy[920], dummy[921], dummy[922], dummy[923], dummy[924], dummy[925], dummy[926], dummy[927], dummy[928], dummy[929], dummy[930], dummy[931], dummy[932], dummy[933], dummy[934], dummy[935], dummy[936], dummy[937], dummy[938], dummy[939], dummy[940], dummy[941], dummy[942], dummy[943], dummy[944], dummy[945], dummy[946], dummy[947], dummy[948], dummy[949], dummy[950], dummy[951], dummy[952], dummy[953], dummy[954], dummy[955], dummy[956], dummy[957], dummy[958], dummy[959], dummy[960], dummy[961], dummy[962], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f963( dummy[963], vec_63_bits[19], vec_63_bits[18] );
    foobar f964( dummy[964], vec_63_bits[20], vec_63_bits[18] );
    foobar f965( dummy[965], vec_63_bits[21], vec_63_bits[18] );
    foobar f966( dummy[966], vec_63_bits[22], vec_63_bits[18] );
    foobar f967( dummy[967], vec_63_bits[23], vec_63_bits[18] );
    foobar f968( dummy[968], vec_63_bits[24], vec_63_bits[18] );
    foobar f969( dummy[969], vec_63_bits[25], vec_63_bits[18] );
    foobar f970( dummy[970], vec_63_bits[26], vec_63_bits[18] );
    foobar f971( dummy[971], vec_63_bits[27], vec_63_bits[18] );
    foobar f972( dummy[972], vec_63_bits[28], vec_63_bits[18] );
    foobar f973( dummy[973], vec_63_bits[29], vec_63_bits[18] );
    foobar f974( dummy[974], vec_63_bits[30], vec_63_bits[18] );
    foobar f975( dummy[975], vec_63_bits[31], vec_63_bits[18] );
    foobar f976( dummy[976], vec_63_bits[32], vec_63_bits[18] );
    foobar f977( dummy[977], vec_63_bits[33], vec_63_bits[18] );
    foobar f978( dummy[978], vec_63_bits[34], vec_63_bits[18] );
    foobar f979( dummy[979], vec_63_bits[35], vec_63_bits[18] );
    foobar f980( dummy[980], vec_63_bits[36], vec_63_bits[18] );
    foobar f981( dummy[981], vec_63_bits[37], vec_63_bits[18] );
    foobar f982( dummy[982], vec_63_bits[38], vec_63_bits[18] );
    foobar f983( dummy[983], vec_63_bits[39], vec_63_bits[18] );
    foobar f984( dummy[984], vec_63_bits[40], vec_63_bits[18] );
    foobar f985( dummy[985], vec_63_bits[41], vec_63_bits[18] );
    foobar f986( dummy[986], vec_63_bits[42], vec_63_bits[18] );
    foobar f987( dummy[987], vec_63_bits[43], vec_63_bits[18] );
    foobar f988( dummy[988], vec_63_bits[44], vec_63_bits[18] );
    foobar f989( dummy[989], vec_63_bits[45], vec_63_bits[18] );
    foobar f990( dummy[990], vec_63_bits[46], vec_63_bits[18] );
    foobar f991( dummy[991], vec_63_bits[47], vec_63_bits[18] );
    foobar f992( dummy[992], vec_63_bits[48], vec_63_bits[18] );
    foobar f993( dummy[993], vec_63_bits[49], vec_63_bits[18] );
    foobar f994( dummy[994], vec_63_bits[50], vec_63_bits[18] );
    foobar f995( dummy[995], vec_63_bits[51], vec_63_bits[18] );
    foobar f996( dummy[996], vec_63_bits[52], vec_63_bits[18] );
    foobar f997( dummy[997], vec_63_bits[53], vec_63_bits[18] );
    foobar f998( dummy[998], vec_63_bits[54], vec_63_bits[18] );
    foobar f999( dummy[999], vec_63_bits[55], vec_63_bits[18] );
    foobar f1000( dummy[1000], vec_63_bits[56], vec_63_bits[18] );
    foobar f1001( dummy[1001], vec_63_bits[57], vec_63_bits[18] );
    foobar f1002( dummy[1002], vec_63_bits[58], vec_63_bits[18] );
    foobar f1003( dummy[1003], vec_63_bits[59], vec_63_bits[18] );
    foobar f1004( dummy[1004], vec_63_bits[60], vec_63_bits[18] );
    foobar f1005( dummy[1005], vec_63_bits[61], vec_63_bits[18] );
    foobar f1006( dummy[1006], vec_63_bits[62], vec_63_bits[18] );
    AN64   an18( o[18], {dummy[963], dummy[964], dummy[965], dummy[966], dummy[967], dummy[968], dummy[969], dummy[970], dummy[971], dummy[972], dummy[973], dummy[974], dummy[975], dummy[976], dummy[977], dummy[978], dummy[979], dummy[980], dummy[981], dummy[982], dummy[983], dummy[984], dummy[985], dummy[986], dummy[987], dummy[988], dummy[989], dummy[990], dummy[991], dummy[992], dummy[993], dummy[994], dummy[995], dummy[996], dummy[997], dummy[998], dummy[999], dummy[1000], dummy[1001], dummy[1002], dummy[1003], dummy[1004], dummy[1005], dummy[1006], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1007( dummy[1007], vec_63_bits[20], vec_63_bits[19] );
    foobar f1008( dummy[1008], vec_63_bits[21], vec_63_bits[19] );
    foobar f1009( dummy[1009], vec_63_bits[22], vec_63_bits[19] );
    foobar f1010( dummy[1010], vec_63_bits[23], vec_63_bits[19] );
    foobar f1011( dummy[1011], vec_63_bits[24], vec_63_bits[19] );
    foobar f1012( dummy[1012], vec_63_bits[25], vec_63_bits[19] );
    foobar f1013( dummy[1013], vec_63_bits[26], vec_63_bits[19] );
    foobar f1014( dummy[1014], vec_63_bits[27], vec_63_bits[19] );
    foobar f1015( dummy[1015], vec_63_bits[28], vec_63_bits[19] );
    foobar f1016( dummy[1016], vec_63_bits[29], vec_63_bits[19] );
    foobar f1017( dummy[1017], vec_63_bits[30], vec_63_bits[19] );
    foobar f1018( dummy[1018], vec_63_bits[31], vec_63_bits[19] );
    foobar f1019( dummy[1019], vec_63_bits[32], vec_63_bits[19] );
    foobar f1020( dummy[1020], vec_63_bits[33], vec_63_bits[19] );
    foobar f1021( dummy[1021], vec_63_bits[34], vec_63_bits[19] );
    foobar f1022( dummy[1022], vec_63_bits[35], vec_63_bits[19] );
    foobar f1023( dummy[1023], vec_63_bits[36], vec_63_bits[19] );
    foobar f1024( dummy[1024], vec_63_bits[37], vec_63_bits[19] );
    foobar f1025( dummy[1025], vec_63_bits[38], vec_63_bits[19] );
    foobar f1026( dummy[1026], vec_63_bits[39], vec_63_bits[19] );
    foobar f1027( dummy[1027], vec_63_bits[40], vec_63_bits[19] );
    foobar f1028( dummy[1028], vec_63_bits[41], vec_63_bits[19] );
    foobar f1029( dummy[1029], vec_63_bits[42], vec_63_bits[19] );
    foobar f1030( dummy[1030], vec_63_bits[43], vec_63_bits[19] );
    foobar f1031( dummy[1031], vec_63_bits[44], vec_63_bits[19] );
    foobar f1032( dummy[1032], vec_63_bits[45], vec_63_bits[19] );
    foobar f1033( dummy[1033], vec_63_bits[46], vec_63_bits[19] );
    foobar f1034( dummy[1034], vec_63_bits[47], vec_63_bits[19] );
    foobar f1035( dummy[1035], vec_63_bits[48], vec_63_bits[19] );
    foobar f1036( dummy[1036], vec_63_bits[49], vec_63_bits[19] );
    foobar f1037( dummy[1037], vec_63_bits[50], vec_63_bits[19] );
    foobar f1038( dummy[1038], vec_63_bits[51], vec_63_bits[19] );
    foobar f1039( dummy[1039], vec_63_bits[52], vec_63_bits[19] );
    foobar f1040( dummy[1040], vec_63_bits[53], vec_63_bits[19] );
    foobar f1041( dummy[1041], vec_63_bits[54], vec_63_bits[19] );
    foobar f1042( dummy[1042], vec_63_bits[55], vec_63_bits[19] );
    foobar f1043( dummy[1043], vec_63_bits[56], vec_63_bits[19] );
    foobar f1044( dummy[1044], vec_63_bits[57], vec_63_bits[19] );
    foobar f1045( dummy[1045], vec_63_bits[58], vec_63_bits[19] );
    foobar f1046( dummy[1046], vec_63_bits[59], vec_63_bits[19] );
    foobar f1047( dummy[1047], vec_63_bits[60], vec_63_bits[19] );
    foobar f1048( dummy[1048], vec_63_bits[61], vec_63_bits[19] );
    foobar f1049( dummy[1049], vec_63_bits[62], vec_63_bits[19] );
    AN64   an19( o[19], {dummy[1007], dummy[1008], dummy[1009], dummy[1010], dummy[1011], dummy[1012], dummy[1013], dummy[1014], dummy[1015], dummy[1016], dummy[1017], dummy[1018], dummy[1019], dummy[1020], dummy[1021], dummy[1022], dummy[1023], dummy[1024], dummy[1025], dummy[1026], dummy[1027], dummy[1028], dummy[1029], dummy[1030], dummy[1031], dummy[1032], dummy[1033], dummy[1034], dummy[1035], dummy[1036], dummy[1037], dummy[1038], dummy[1039], dummy[1040], dummy[1041], dummy[1042], dummy[1043], dummy[1044], dummy[1045], dummy[1046], dummy[1047], dummy[1048], dummy[1049], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1050( dummy[1050], vec_63_bits[21], vec_63_bits[20] );
    foobar f1051( dummy[1051], vec_63_bits[22], vec_63_bits[20] );
    foobar f1052( dummy[1052], vec_63_bits[23], vec_63_bits[20] );
    foobar f1053( dummy[1053], vec_63_bits[24], vec_63_bits[20] );
    foobar f1054( dummy[1054], vec_63_bits[25], vec_63_bits[20] );
    foobar f1055( dummy[1055], vec_63_bits[26], vec_63_bits[20] );
    foobar f1056( dummy[1056], vec_63_bits[27], vec_63_bits[20] );
    foobar f1057( dummy[1057], vec_63_bits[28], vec_63_bits[20] );
    foobar f1058( dummy[1058], vec_63_bits[29], vec_63_bits[20] );
    foobar f1059( dummy[1059], vec_63_bits[30], vec_63_bits[20] );
    foobar f1060( dummy[1060], vec_63_bits[31], vec_63_bits[20] );
    foobar f1061( dummy[1061], vec_63_bits[32], vec_63_bits[20] );
    foobar f1062( dummy[1062], vec_63_bits[33], vec_63_bits[20] );
    foobar f1063( dummy[1063], vec_63_bits[34], vec_63_bits[20] );
    foobar f1064( dummy[1064], vec_63_bits[35], vec_63_bits[20] );
    foobar f1065( dummy[1065], vec_63_bits[36], vec_63_bits[20] );
    foobar f1066( dummy[1066], vec_63_bits[37], vec_63_bits[20] );
    foobar f1067( dummy[1067], vec_63_bits[38], vec_63_bits[20] );
    foobar f1068( dummy[1068], vec_63_bits[39], vec_63_bits[20] );
    foobar f1069( dummy[1069], vec_63_bits[40], vec_63_bits[20] );
    foobar f1070( dummy[1070], vec_63_bits[41], vec_63_bits[20] );
    foobar f1071( dummy[1071], vec_63_bits[42], vec_63_bits[20] );
    foobar f1072( dummy[1072], vec_63_bits[43], vec_63_bits[20] );
    foobar f1073( dummy[1073], vec_63_bits[44], vec_63_bits[20] );
    foobar f1074( dummy[1074], vec_63_bits[45], vec_63_bits[20] );
    foobar f1075( dummy[1075], vec_63_bits[46], vec_63_bits[20] );
    foobar f1076( dummy[1076], vec_63_bits[47], vec_63_bits[20] );
    foobar f1077( dummy[1077], vec_63_bits[48], vec_63_bits[20] );
    foobar f1078( dummy[1078], vec_63_bits[49], vec_63_bits[20] );
    foobar f1079( dummy[1079], vec_63_bits[50], vec_63_bits[20] );
    foobar f1080( dummy[1080], vec_63_bits[51], vec_63_bits[20] );
    foobar f1081( dummy[1081], vec_63_bits[52], vec_63_bits[20] );
    foobar f1082( dummy[1082], vec_63_bits[53], vec_63_bits[20] );
    foobar f1083( dummy[1083], vec_63_bits[54], vec_63_bits[20] );
    foobar f1084( dummy[1084], vec_63_bits[55], vec_63_bits[20] );
    foobar f1085( dummy[1085], vec_63_bits[56], vec_63_bits[20] );
    foobar f1086( dummy[1086], vec_63_bits[57], vec_63_bits[20] );
    foobar f1087( dummy[1087], vec_63_bits[58], vec_63_bits[20] );
    foobar f1088( dummy[1088], vec_63_bits[59], vec_63_bits[20] );
    foobar f1089( dummy[1089], vec_63_bits[60], vec_63_bits[20] );
    foobar f1090( dummy[1090], vec_63_bits[61], vec_63_bits[20] );
    foobar f1091( dummy[1091], vec_63_bits[62], vec_63_bits[20] );
    AN64   an20( o[20], {dummy[1050], dummy[1051], dummy[1052], dummy[1053], dummy[1054], dummy[1055], dummy[1056], dummy[1057], dummy[1058], dummy[1059], dummy[1060], dummy[1061], dummy[1062], dummy[1063], dummy[1064], dummy[1065], dummy[1066], dummy[1067], dummy[1068], dummy[1069], dummy[1070], dummy[1071], dummy[1072], dummy[1073], dummy[1074], dummy[1075], dummy[1076], dummy[1077], dummy[1078], dummy[1079], dummy[1080], dummy[1081], dummy[1082], dummy[1083], dummy[1084], dummy[1085], dummy[1086], dummy[1087], dummy[1088], dummy[1089], dummy[1090], dummy[1091], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1092( dummy[1092], vec_63_bits[22], vec_63_bits[21] );
    foobar f1093( dummy[1093], vec_63_bits[23], vec_63_bits[21] );
    foobar f1094( dummy[1094], vec_63_bits[24], vec_63_bits[21] );
    foobar f1095( dummy[1095], vec_63_bits[25], vec_63_bits[21] );
    foobar f1096( dummy[1096], vec_63_bits[26], vec_63_bits[21] );
    foobar f1097( dummy[1097], vec_63_bits[27], vec_63_bits[21] );
    foobar f1098( dummy[1098], vec_63_bits[28], vec_63_bits[21] );
    foobar f1099( dummy[1099], vec_63_bits[29], vec_63_bits[21] );
    foobar f1100( dummy[1100], vec_63_bits[30], vec_63_bits[21] );
    foobar f1101( dummy[1101], vec_63_bits[31], vec_63_bits[21] );
    foobar f1102( dummy[1102], vec_63_bits[32], vec_63_bits[21] );
    foobar f1103( dummy[1103], vec_63_bits[33], vec_63_bits[21] );
    foobar f1104( dummy[1104], vec_63_bits[34], vec_63_bits[21] );
    foobar f1105( dummy[1105], vec_63_bits[35], vec_63_bits[21] );
    foobar f1106( dummy[1106], vec_63_bits[36], vec_63_bits[21] );
    foobar f1107( dummy[1107], vec_63_bits[37], vec_63_bits[21] );
    foobar f1108( dummy[1108], vec_63_bits[38], vec_63_bits[21] );
    foobar f1109( dummy[1109], vec_63_bits[39], vec_63_bits[21] );
    foobar f1110( dummy[1110], vec_63_bits[40], vec_63_bits[21] );
    foobar f1111( dummy[1111], vec_63_bits[41], vec_63_bits[21] );
    foobar f1112( dummy[1112], vec_63_bits[42], vec_63_bits[21] );
    foobar f1113( dummy[1113], vec_63_bits[43], vec_63_bits[21] );
    foobar f1114( dummy[1114], vec_63_bits[44], vec_63_bits[21] );
    foobar f1115( dummy[1115], vec_63_bits[45], vec_63_bits[21] );
    foobar f1116( dummy[1116], vec_63_bits[46], vec_63_bits[21] );
    foobar f1117( dummy[1117], vec_63_bits[47], vec_63_bits[21] );
    foobar f1118( dummy[1118], vec_63_bits[48], vec_63_bits[21] );
    foobar f1119( dummy[1119], vec_63_bits[49], vec_63_bits[21] );
    foobar f1120( dummy[1120], vec_63_bits[50], vec_63_bits[21] );
    foobar f1121( dummy[1121], vec_63_bits[51], vec_63_bits[21] );
    foobar f1122( dummy[1122], vec_63_bits[52], vec_63_bits[21] );
    foobar f1123( dummy[1123], vec_63_bits[53], vec_63_bits[21] );
    foobar f1124( dummy[1124], vec_63_bits[54], vec_63_bits[21] );
    foobar f1125( dummy[1125], vec_63_bits[55], vec_63_bits[21] );
    foobar f1126( dummy[1126], vec_63_bits[56], vec_63_bits[21] );
    foobar f1127( dummy[1127], vec_63_bits[57], vec_63_bits[21] );
    foobar f1128( dummy[1128], vec_63_bits[58], vec_63_bits[21] );
    foobar f1129( dummy[1129], vec_63_bits[59], vec_63_bits[21] );
    foobar f1130( dummy[1130], vec_63_bits[60], vec_63_bits[21] );
    foobar f1131( dummy[1131], vec_63_bits[61], vec_63_bits[21] );
    foobar f1132( dummy[1132], vec_63_bits[62], vec_63_bits[21] );
    AN64   an21( o[21], {dummy[1092], dummy[1093], dummy[1094], dummy[1095], dummy[1096], dummy[1097], dummy[1098], dummy[1099], dummy[1100], dummy[1101], dummy[1102], dummy[1103], dummy[1104], dummy[1105], dummy[1106], dummy[1107], dummy[1108], dummy[1109], dummy[1110], dummy[1111], dummy[1112], dummy[1113], dummy[1114], dummy[1115], dummy[1116], dummy[1117], dummy[1118], dummy[1119], dummy[1120], dummy[1121], dummy[1122], dummy[1123], dummy[1124], dummy[1125], dummy[1126], dummy[1127], dummy[1128], dummy[1129], dummy[1130], dummy[1131], dummy[1132], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1133( dummy[1133], vec_63_bits[23], vec_63_bits[22] );
    foobar f1134( dummy[1134], vec_63_bits[24], vec_63_bits[22] );
    foobar f1135( dummy[1135], vec_63_bits[25], vec_63_bits[22] );
    foobar f1136( dummy[1136], vec_63_bits[26], vec_63_bits[22] );
    foobar f1137( dummy[1137], vec_63_bits[27], vec_63_bits[22] );
    foobar f1138( dummy[1138], vec_63_bits[28], vec_63_bits[22] );
    foobar f1139( dummy[1139], vec_63_bits[29], vec_63_bits[22] );
    foobar f1140( dummy[1140], vec_63_bits[30], vec_63_bits[22] );
    foobar f1141( dummy[1141], vec_63_bits[31], vec_63_bits[22] );
    foobar f1142( dummy[1142], vec_63_bits[32], vec_63_bits[22] );
    foobar f1143( dummy[1143], vec_63_bits[33], vec_63_bits[22] );
    foobar f1144( dummy[1144], vec_63_bits[34], vec_63_bits[22] );
    foobar f1145( dummy[1145], vec_63_bits[35], vec_63_bits[22] );
    foobar f1146( dummy[1146], vec_63_bits[36], vec_63_bits[22] );
    foobar f1147( dummy[1147], vec_63_bits[37], vec_63_bits[22] );
    foobar f1148( dummy[1148], vec_63_bits[38], vec_63_bits[22] );
    foobar f1149( dummy[1149], vec_63_bits[39], vec_63_bits[22] );
    foobar f1150( dummy[1150], vec_63_bits[40], vec_63_bits[22] );
    foobar f1151( dummy[1151], vec_63_bits[41], vec_63_bits[22] );
    foobar f1152( dummy[1152], vec_63_bits[42], vec_63_bits[22] );
    foobar f1153( dummy[1153], vec_63_bits[43], vec_63_bits[22] );
    foobar f1154( dummy[1154], vec_63_bits[44], vec_63_bits[22] );
    foobar f1155( dummy[1155], vec_63_bits[45], vec_63_bits[22] );
    foobar f1156( dummy[1156], vec_63_bits[46], vec_63_bits[22] );
    foobar f1157( dummy[1157], vec_63_bits[47], vec_63_bits[22] );
    foobar f1158( dummy[1158], vec_63_bits[48], vec_63_bits[22] );
    foobar f1159( dummy[1159], vec_63_bits[49], vec_63_bits[22] );
    foobar f1160( dummy[1160], vec_63_bits[50], vec_63_bits[22] );
    foobar f1161( dummy[1161], vec_63_bits[51], vec_63_bits[22] );
    foobar f1162( dummy[1162], vec_63_bits[52], vec_63_bits[22] );
    foobar f1163( dummy[1163], vec_63_bits[53], vec_63_bits[22] );
    foobar f1164( dummy[1164], vec_63_bits[54], vec_63_bits[22] );
    foobar f1165( dummy[1165], vec_63_bits[55], vec_63_bits[22] );
    foobar f1166( dummy[1166], vec_63_bits[56], vec_63_bits[22] );
    foobar f1167( dummy[1167], vec_63_bits[57], vec_63_bits[22] );
    foobar f1168( dummy[1168], vec_63_bits[58], vec_63_bits[22] );
    foobar f1169( dummy[1169], vec_63_bits[59], vec_63_bits[22] );
    foobar f1170( dummy[1170], vec_63_bits[60], vec_63_bits[22] );
    foobar f1171( dummy[1171], vec_63_bits[61], vec_63_bits[22] );
    foobar f1172( dummy[1172], vec_63_bits[62], vec_63_bits[22] );
    AN64   an22( o[22], {dummy[1133], dummy[1134], dummy[1135], dummy[1136], dummy[1137], dummy[1138], dummy[1139], dummy[1140], dummy[1141], dummy[1142], dummy[1143], dummy[1144], dummy[1145], dummy[1146], dummy[1147], dummy[1148], dummy[1149], dummy[1150], dummy[1151], dummy[1152], dummy[1153], dummy[1154], dummy[1155], dummy[1156], dummy[1157], dummy[1158], dummy[1159], dummy[1160], dummy[1161], dummy[1162], dummy[1163], dummy[1164], dummy[1165], dummy[1166], dummy[1167], dummy[1168], dummy[1169], dummy[1170], dummy[1171], dummy[1172], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1173( dummy[1173], vec_63_bits[24], vec_63_bits[23] );
    foobar f1174( dummy[1174], vec_63_bits[25], vec_63_bits[23] );
    foobar f1175( dummy[1175], vec_63_bits[26], vec_63_bits[23] );
    foobar f1176( dummy[1176], vec_63_bits[27], vec_63_bits[23] );
    foobar f1177( dummy[1177], vec_63_bits[28], vec_63_bits[23] );
    foobar f1178( dummy[1178], vec_63_bits[29], vec_63_bits[23] );
    foobar f1179( dummy[1179], vec_63_bits[30], vec_63_bits[23] );
    foobar f1180( dummy[1180], vec_63_bits[31], vec_63_bits[23] );
    foobar f1181( dummy[1181], vec_63_bits[32], vec_63_bits[23] );
    foobar f1182( dummy[1182], vec_63_bits[33], vec_63_bits[23] );
    foobar f1183( dummy[1183], vec_63_bits[34], vec_63_bits[23] );
    foobar f1184( dummy[1184], vec_63_bits[35], vec_63_bits[23] );
    foobar f1185( dummy[1185], vec_63_bits[36], vec_63_bits[23] );
    foobar f1186( dummy[1186], vec_63_bits[37], vec_63_bits[23] );
    foobar f1187( dummy[1187], vec_63_bits[38], vec_63_bits[23] );
    foobar f1188( dummy[1188], vec_63_bits[39], vec_63_bits[23] );
    foobar f1189( dummy[1189], vec_63_bits[40], vec_63_bits[23] );
    foobar f1190( dummy[1190], vec_63_bits[41], vec_63_bits[23] );
    foobar f1191( dummy[1191], vec_63_bits[42], vec_63_bits[23] );
    foobar f1192( dummy[1192], vec_63_bits[43], vec_63_bits[23] );
    foobar f1193( dummy[1193], vec_63_bits[44], vec_63_bits[23] );
    foobar f1194( dummy[1194], vec_63_bits[45], vec_63_bits[23] );
    foobar f1195( dummy[1195], vec_63_bits[46], vec_63_bits[23] );
    foobar f1196( dummy[1196], vec_63_bits[47], vec_63_bits[23] );
    foobar f1197( dummy[1197], vec_63_bits[48], vec_63_bits[23] );
    foobar f1198( dummy[1198], vec_63_bits[49], vec_63_bits[23] );
    foobar f1199( dummy[1199], vec_63_bits[50], vec_63_bits[23] );
    foobar f1200( dummy[1200], vec_63_bits[51], vec_63_bits[23] );
    foobar f1201( dummy[1201], vec_63_bits[52], vec_63_bits[23] );
    foobar f1202( dummy[1202], vec_63_bits[53], vec_63_bits[23] );
    foobar f1203( dummy[1203], vec_63_bits[54], vec_63_bits[23] );
    foobar f1204( dummy[1204], vec_63_bits[55], vec_63_bits[23] );
    foobar f1205( dummy[1205], vec_63_bits[56], vec_63_bits[23] );
    foobar f1206( dummy[1206], vec_63_bits[57], vec_63_bits[23] );
    foobar f1207( dummy[1207], vec_63_bits[58], vec_63_bits[23] );
    foobar f1208( dummy[1208], vec_63_bits[59], vec_63_bits[23] );
    foobar f1209( dummy[1209], vec_63_bits[60], vec_63_bits[23] );
    foobar f1210( dummy[1210], vec_63_bits[61], vec_63_bits[23] );
    foobar f1211( dummy[1211], vec_63_bits[62], vec_63_bits[23] );
    AN64   an23( o[23], {dummy[1173], dummy[1174], dummy[1175], dummy[1176], dummy[1177], dummy[1178], dummy[1179], dummy[1180], dummy[1181], dummy[1182], dummy[1183], dummy[1184], dummy[1185], dummy[1186], dummy[1187], dummy[1188], dummy[1189], dummy[1190], dummy[1191], dummy[1192], dummy[1193], dummy[1194], dummy[1195], dummy[1196], dummy[1197], dummy[1198], dummy[1199], dummy[1200], dummy[1201], dummy[1202], dummy[1203], dummy[1204], dummy[1205], dummy[1206], dummy[1207], dummy[1208], dummy[1209], dummy[1210], dummy[1211], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1212( dummy[1212], vec_63_bits[25], vec_63_bits[24] );
    foobar f1213( dummy[1213], vec_63_bits[26], vec_63_bits[24] );
    foobar f1214( dummy[1214], vec_63_bits[27], vec_63_bits[24] );
    foobar f1215( dummy[1215], vec_63_bits[28], vec_63_bits[24] );
    foobar f1216( dummy[1216], vec_63_bits[29], vec_63_bits[24] );
    foobar f1217( dummy[1217], vec_63_bits[30], vec_63_bits[24] );
    foobar f1218( dummy[1218], vec_63_bits[31], vec_63_bits[24] );
    foobar f1219( dummy[1219], vec_63_bits[32], vec_63_bits[24] );
    foobar f1220( dummy[1220], vec_63_bits[33], vec_63_bits[24] );
    foobar f1221( dummy[1221], vec_63_bits[34], vec_63_bits[24] );
    foobar f1222( dummy[1222], vec_63_bits[35], vec_63_bits[24] );
    foobar f1223( dummy[1223], vec_63_bits[36], vec_63_bits[24] );
    foobar f1224( dummy[1224], vec_63_bits[37], vec_63_bits[24] );
    foobar f1225( dummy[1225], vec_63_bits[38], vec_63_bits[24] );
    foobar f1226( dummy[1226], vec_63_bits[39], vec_63_bits[24] );
    foobar f1227( dummy[1227], vec_63_bits[40], vec_63_bits[24] );
    foobar f1228( dummy[1228], vec_63_bits[41], vec_63_bits[24] );
    foobar f1229( dummy[1229], vec_63_bits[42], vec_63_bits[24] );
    foobar f1230( dummy[1230], vec_63_bits[43], vec_63_bits[24] );
    foobar f1231( dummy[1231], vec_63_bits[44], vec_63_bits[24] );
    foobar f1232( dummy[1232], vec_63_bits[45], vec_63_bits[24] );
    foobar f1233( dummy[1233], vec_63_bits[46], vec_63_bits[24] );
    foobar f1234( dummy[1234], vec_63_bits[47], vec_63_bits[24] );
    foobar f1235( dummy[1235], vec_63_bits[48], vec_63_bits[24] );
    foobar f1236( dummy[1236], vec_63_bits[49], vec_63_bits[24] );
    foobar f1237( dummy[1237], vec_63_bits[50], vec_63_bits[24] );
    foobar f1238( dummy[1238], vec_63_bits[51], vec_63_bits[24] );
    foobar f1239( dummy[1239], vec_63_bits[52], vec_63_bits[24] );
    foobar f1240( dummy[1240], vec_63_bits[53], vec_63_bits[24] );
    foobar f1241( dummy[1241], vec_63_bits[54], vec_63_bits[24] );
    foobar f1242( dummy[1242], vec_63_bits[55], vec_63_bits[24] );
    foobar f1243( dummy[1243], vec_63_bits[56], vec_63_bits[24] );
    foobar f1244( dummy[1244], vec_63_bits[57], vec_63_bits[24] );
    foobar f1245( dummy[1245], vec_63_bits[58], vec_63_bits[24] );
    foobar f1246( dummy[1246], vec_63_bits[59], vec_63_bits[24] );
    foobar f1247( dummy[1247], vec_63_bits[60], vec_63_bits[24] );
    foobar f1248( dummy[1248], vec_63_bits[61], vec_63_bits[24] );
    foobar f1249( dummy[1249], vec_63_bits[62], vec_63_bits[24] );
    AN64   an24( o[24], {dummy[1212], dummy[1213], dummy[1214], dummy[1215], dummy[1216], dummy[1217], dummy[1218], dummy[1219], dummy[1220], dummy[1221], dummy[1222], dummy[1223], dummy[1224], dummy[1225], dummy[1226], dummy[1227], dummy[1228], dummy[1229], dummy[1230], dummy[1231], dummy[1232], dummy[1233], dummy[1234], dummy[1235], dummy[1236], dummy[1237], dummy[1238], dummy[1239], dummy[1240], dummy[1241], dummy[1242], dummy[1243], dummy[1244], dummy[1245], dummy[1246], dummy[1247], dummy[1248], dummy[1249], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1250( dummy[1250], vec_63_bits[26], vec_63_bits[25] );
    foobar f1251( dummy[1251], vec_63_bits[27], vec_63_bits[25] );
    foobar f1252( dummy[1252], vec_63_bits[28], vec_63_bits[25] );
    foobar f1253( dummy[1253], vec_63_bits[29], vec_63_bits[25] );
    foobar f1254( dummy[1254], vec_63_bits[30], vec_63_bits[25] );
    foobar f1255( dummy[1255], vec_63_bits[31], vec_63_bits[25] );
    foobar f1256( dummy[1256], vec_63_bits[32], vec_63_bits[25] );
    foobar f1257( dummy[1257], vec_63_bits[33], vec_63_bits[25] );
    foobar f1258( dummy[1258], vec_63_bits[34], vec_63_bits[25] );
    foobar f1259( dummy[1259], vec_63_bits[35], vec_63_bits[25] );
    foobar f1260( dummy[1260], vec_63_bits[36], vec_63_bits[25] );
    foobar f1261( dummy[1261], vec_63_bits[37], vec_63_bits[25] );
    foobar f1262( dummy[1262], vec_63_bits[38], vec_63_bits[25] );
    foobar f1263( dummy[1263], vec_63_bits[39], vec_63_bits[25] );
    foobar f1264( dummy[1264], vec_63_bits[40], vec_63_bits[25] );
    foobar f1265( dummy[1265], vec_63_bits[41], vec_63_bits[25] );
    foobar f1266( dummy[1266], vec_63_bits[42], vec_63_bits[25] );
    foobar f1267( dummy[1267], vec_63_bits[43], vec_63_bits[25] );
    foobar f1268( dummy[1268], vec_63_bits[44], vec_63_bits[25] );
    foobar f1269( dummy[1269], vec_63_bits[45], vec_63_bits[25] );
    foobar f1270( dummy[1270], vec_63_bits[46], vec_63_bits[25] );
    foobar f1271( dummy[1271], vec_63_bits[47], vec_63_bits[25] );
    foobar f1272( dummy[1272], vec_63_bits[48], vec_63_bits[25] );
    foobar f1273( dummy[1273], vec_63_bits[49], vec_63_bits[25] );
    foobar f1274( dummy[1274], vec_63_bits[50], vec_63_bits[25] );
    foobar f1275( dummy[1275], vec_63_bits[51], vec_63_bits[25] );
    foobar f1276( dummy[1276], vec_63_bits[52], vec_63_bits[25] );
    foobar f1277( dummy[1277], vec_63_bits[53], vec_63_bits[25] );
    foobar f1278( dummy[1278], vec_63_bits[54], vec_63_bits[25] );
    foobar f1279( dummy[1279], vec_63_bits[55], vec_63_bits[25] );
    foobar f1280( dummy[1280], vec_63_bits[56], vec_63_bits[25] );
    foobar f1281( dummy[1281], vec_63_bits[57], vec_63_bits[25] );
    foobar f1282( dummy[1282], vec_63_bits[58], vec_63_bits[25] );
    foobar f1283( dummy[1283], vec_63_bits[59], vec_63_bits[25] );
    foobar f1284( dummy[1284], vec_63_bits[60], vec_63_bits[25] );
    foobar f1285( dummy[1285], vec_63_bits[61], vec_63_bits[25] );
    foobar f1286( dummy[1286], vec_63_bits[62], vec_63_bits[25] );
    AN64   an25( o[25], {dummy[1250], dummy[1251], dummy[1252], dummy[1253], dummy[1254], dummy[1255], dummy[1256], dummy[1257], dummy[1258], dummy[1259], dummy[1260], dummy[1261], dummy[1262], dummy[1263], dummy[1264], dummy[1265], dummy[1266], dummy[1267], dummy[1268], dummy[1269], dummy[1270], dummy[1271], dummy[1272], dummy[1273], dummy[1274], dummy[1275], dummy[1276], dummy[1277], dummy[1278], dummy[1279], dummy[1280], dummy[1281], dummy[1282], dummy[1283], dummy[1284], dummy[1285], dummy[1286], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1287( dummy[1287], vec_63_bits[27], vec_63_bits[26] );
    foobar f1288( dummy[1288], vec_63_bits[28], vec_63_bits[26] );
    foobar f1289( dummy[1289], vec_63_bits[29], vec_63_bits[26] );
    foobar f1290( dummy[1290], vec_63_bits[30], vec_63_bits[26] );
    foobar f1291( dummy[1291], vec_63_bits[31], vec_63_bits[26] );
    foobar f1292( dummy[1292], vec_63_bits[32], vec_63_bits[26] );
    foobar f1293( dummy[1293], vec_63_bits[33], vec_63_bits[26] );
    foobar f1294( dummy[1294], vec_63_bits[34], vec_63_bits[26] );
    foobar f1295( dummy[1295], vec_63_bits[35], vec_63_bits[26] );
    foobar f1296( dummy[1296], vec_63_bits[36], vec_63_bits[26] );
    foobar f1297( dummy[1297], vec_63_bits[37], vec_63_bits[26] );
    foobar f1298( dummy[1298], vec_63_bits[38], vec_63_bits[26] );
    foobar f1299( dummy[1299], vec_63_bits[39], vec_63_bits[26] );
    foobar f1300( dummy[1300], vec_63_bits[40], vec_63_bits[26] );
    foobar f1301( dummy[1301], vec_63_bits[41], vec_63_bits[26] );
    foobar f1302( dummy[1302], vec_63_bits[42], vec_63_bits[26] );
    foobar f1303( dummy[1303], vec_63_bits[43], vec_63_bits[26] );
    foobar f1304( dummy[1304], vec_63_bits[44], vec_63_bits[26] );
    foobar f1305( dummy[1305], vec_63_bits[45], vec_63_bits[26] );
    foobar f1306( dummy[1306], vec_63_bits[46], vec_63_bits[26] );
    foobar f1307( dummy[1307], vec_63_bits[47], vec_63_bits[26] );
    foobar f1308( dummy[1308], vec_63_bits[48], vec_63_bits[26] );
    foobar f1309( dummy[1309], vec_63_bits[49], vec_63_bits[26] );
    foobar f1310( dummy[1310], vec_63_bits[50], vec_63_bits[26] );
    foobar f1311( dummy[1311], vec_63_bits[51], vec_63_bits[26] );
    foobar f1312( dummy[1312], vec_63_bits[52], vec_63_bits[26] );
    foobar f1313( dummy[1313], vec_63_bits[53], vec_63_bits[26] );
    foobar f1314( dummy[1314], vec_63_bits[54], vec_63_bits[26] );
    foobar f1315( dummy[1315], vec_63_bits[55], vec_63_bits[26] );
    foobar f1316( dummy[1316], vec_63_bits[56], vec_63_bits[26] );
    foobar f1317( dummy[1317], vec_63_bits[57], vec_63_bits[26] );
    foobar f1318( dummy[1318], vec_63_bits[58], vec_63_bits[26] );
    foobar f1319( dummy[1319], vec_63_bits[59], vec_63_bits[26] );
    foobar f1320( dummy[1320], vec_63_bits[60], vec_63_bits[26] );
    foobar f1321( dummy[1321], vec_63_bits[61], vec_63_bits[26] );
    foobar f1322( dummy[1322], vec_63_bits[62], vec_63_bits[26] );
    AN64   an26( o[26], {dummy[1287], dummy[1288], dummy[1289], dummy[1290], dummy[1291], dummy[1292], dummy[1293], dummy[1294], dummy[1295], dummy[1296], dummy[1297], dummy[1298], dummy[1299], dummy[1300], dummy[1301], dummy[1302], dummy[1303], dummy[1304], dummy[1305], dummy[1306], dummy[1307], dummy[1308], dummy[1309], dummy[1310], dummy[1311], dummy[1312], dummy[1313], dummy[1314], dummy[1315], dummy[1316], dummy[1317], dummy[1318], dummy[1319], dummy[1320], dummy[1321], dummy[1322], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1323( dummy[1323], vec_63_bits[28], vec_63_bits[27] );
    foobar f1324( dummy[1324], vec_63_bits[29], vec_63_bits[27] );
    foobar f1325( dummy[1325], vec_63_bits[30], vec_63_bits[27] );
    foobar f1326( dummy[1326], vec_63_bits[31], vec_63_bits[27] );
    foobar f1327( dummy[1327], vec_63_bits[32], vec_63_bits[27] );
    foobar f1328( dummy[1328], vec_63_bits[33], vec_63_bits[27] );
    foobar f1329( dummy[1329], vec_63_bits[34], vec_63_bits[27] );
    foobar f1330( dummy[1330], vec_63_bits[35], vec_63_bits[27] );
    foobar f1331( dummy[1331], vec_63_bits[36], vec_63_bits[27] );
    foobar f1332( dummy[1332], vec_63_bits[37], vec_63_bits[27] );
    foobar f1333( dummy[1333], vec_63_bits[38], vec_63_bits[27] );
    foobar f1334( dummy[1334], vec_63_bits[39], vec_63_bits[27] );
    foobar f1335( dummy[1335], vec_63_bits[40], vec_63_bits[27] );
    foobar f1336( dummy[1336], vec_63_bits[41], vec_63_bits[27] );
    foobar f1337( dummy[1337], vec_63_bits[42], vec_63_bits[27] );
    foobar f1338( dummy[1338], vec_63_bits[43], vec_63_bits[27] );
    foobar f1339( dummy[1339], vec_63_bits[44], vec_63_bits[27] );
    foobar f1340( dummy[1340], vec_63_bits[45], vec_63_bits[27] );
    foobar f1341( dummy[1341], vec_63_bits[46], vec_63_bits[27] );
    foobar f1342( dummy[1342], vec_63_bits[47], vec_63_bits[27] );
    foobar f1343( dummy[1343], vec_63_bits[48], vec_63_bits[27] );
    foobar f1344( dummy[1344], vec_63_bits[49], vec_63_bits[27] );
    foobar f1345( dummy[1345], vec_63_bits[50], vec_63_bits[27] );
    foobar f1346( dummy[1346], vec_63_bits[51], vec_63_bits[27] );
    foobar f1347( dummy[1347], vec_63_bits[52], vec_63_bits[27] );
    foobar f1348( dummy[1348], vec_63_bits[53], vec_63_bits[27] );
    foobar f1349( dummy[1349], vec_63_bits[54], vec_63_bits[27] );
    foobar f1350( dummy[1350], vec_63_bits[55], vec_63_bits[27] );
    foobar f1351( dummy[1351], vec_63_bits[56], vec_63_bits[27] );
    foobar f1352( dummy[1352], vec_63_bits[57], vec_63_bits[27] );
    foobar f1353( dummy[1353], vec_63_bits[58], vec_63_bits[27] );
    foobar f1354( dummy[1354], vec_63_bits[59], vec_63_bits[27] );
    foobar f1355( dummy[1355], vec_63_bits[60], vec_63_bits[27] );
    foobar f1356( dummy[1356], vec_63_bits[61], vec_63_bits[27] );
    foobar f1357( dummy[1357], vec_63_bits[62], vec_63_bits[27] );
    AN64   an27( o[27], {dummy[1323], dummy[1324], dummy[1325], dummy[1326], dummy[1327], dummy[1328], dummy[1329], dummy[1330], dummy[1331], dummy[1332], dummy[1333], dummy[1334], dummy[1335], dummy[1336], dummy[1337], dummy[1338], dummy[1339], dummy[1340], dummy[1341], dummy[1342], dummy[1343], dummy[1344], dummy[1345], dummy[1346], dummy[1347], dummy[1348], dummy[1349], dummy[1350], dummy[1351], dummy[1352], dummy[1353], dummy[1354], dummy[1355], dummy[1356], dummy[1357], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1358( dummy[1358], vec_63_bits[29], vec_63_bits[28] );
    foobar f1359( dummy[1359], vec_63_bits[30], vec_63_bits[28] );
    foobar f1360( dummy[1360], vec_63_bits[31], vec_63_bits[28] );
    foobar f1361( dummy[1361], vec_63_bits[32], vec_63_bits[28] );
    foobar f1362( dummy[1362], vec_63_bits[33], vec_63_bits[28] );
    foobar f1363( dummy[1363], vec_63_bits[34], vec_63_bits[28] );
    foobar f1364( dummy[1364], vec_63_bits[35], vec_63_bits[28] );
    foobar f1365( dummy[1365], vec_63_bits[36], vec_63_bits[28] );
    foobar f1366( dummy[1366], vec_63_bits[37], vec_63_bits[28] );
    foobar f1367( dummy[1367], vec_63_bits[38], vec_63_bits[28] );
    foobar f1368( dummy[1368], vec_63_bits[39], vec_63_bits[28] );
    foobar f1369( dummy[1369], vec_63_bits[40], vec_63_bits[28] );
    foobar f1370( dummy[1370], vec_63_bits[41], vec_63_bits[28] );
    foobar f1371( dummy[1371], vec_63_bits[42], vec_63_bits[28] );
    foobar f1372( dummy[1372], vec_63_bits[43], vec_63_bits[28] );
    foobar f1373( dummy[1373], vec_63_bits[44], vec_63_bits[28] );
    foobar f1374( dummy[1374], vec_63_bits[45], vec_63_bits[28] );
    foobar f1375( dummy[1375], vec_63_bits[46], vec_63_bits[28] );
    foobar f1376( dummy[1376], vec_63_bits[47], vec_63_bits[28] );
    foobar f1377( dummy[1377], vec_63_bits[48], vec_63_bits[28] );
    foobar f1378( dummy[1378], vec_63_bits[49], vec_63_bits[28] );
    foobar f1379( dummy[1379], vec_63_bits[50], vec_63_bits[28] );
    foobar f1380( dummy[1380], vec_63_bits[51], vec_63_bits[28] );
    foobar f1381( dummy[1381], vec_63_bits[52], vec_63_bits[28] );
    foobar f1382( dummy[1382], vec_63_bits[53], vec_63_bits[28] );
    foobar f1383( dummy[1383], vec_63_bits[54], vec_63_bits[28] );
    foobar f1384( dummy[1384], vec_63_bits[55], vec_63_bits[28] );
    foobar f1385( dummy[1385], vec_63_bits[56], vec_63_bits[28] );
    foobar f1386( dummy[1386], vec_63_bits[57], vec_63_bits[28] );
    foobar f1387( dummy[1387], vec_63_bits[58], vec_63_bits[28] );
    foobar f1388( dummy[1388], vec_63_bits[59], vec_63_bits[28] );
    foobar f1389( dummy[1389], vec_63_bits[60], vec_63_bits[28] );
    foobar f1390( dummy[1390], vec_63_bits[61], vec_63_bits[28] );
    foobar f1391( dummy[1391], vec_63_bits[62], vec_63_bits[28] );
    AN64   an28( o[28], {dummy[1358], dummy[1359], dummy[1360], dummy[1361], dummy[1362], dummy[1363], dummy[1364], dummy[1365], dummy[1366], dummy[1367], dummy[1368], dummy[1369], dummy[1370], dummy[1371], dummy[1372], dummy[1373], dummy[1374], dummy[1375], dummy[1376], dummy[1377], dummy[1378], dummy[1379], dummy[1380], dummy[1381], dummy[1382], dummy[1383], dummy[1384], dummy[1385], dummy[1386], dummy[1387], dummy[1388], dummy[1389], dummy[1390], dummy[1391], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1392( dummy[1392], vec_63_bits[30], vec_63_bits[29] );
    foobar f1393( dummy[1393], vec_63_bits[31], vec_63_bits[29] );
    foobar f1394( dummy[1394], vec_63_bits[32], vec_63_bits[29] );
    foobar f1395( dummy[1395], vec_63_bits[33], vec_63_bits[29] );
    foobar f1396( dummy[1396], vec_63_bits[34], vec_63_bits[29] );
    foobar f1397( dummy[1397], vec_63_bits[35], vec_63_bits[29] );
    foobar f1398( dummy[1398], vec_63_bits[36], vec_63_bits[29] );
    foobar f1399( dummy[1399], vec_63_bits[37], vec_63_bits[29] );
    foobar f1400( dummy[1400], vec_63_bits[38], vec_63_bits[29] );
    foobar f1401( dummy[1401], vec_63_bits[39], vec_63_bits[29] );
    foobar f1402( dummy[1402], vec_63_bits[40], vec_63_bits[29] );
    foobar f1403( dummy[1403], vec_63_bits[41], vec_63_bits[29] );
    foobar f1404( dummy[1404], vec_63_bits[42], vec_63_bits[29] );
    foobar f1405( dummy[1405], vec_63_bits[43], vec_63_bits[29] );
    foobar f1406( dummy[1406], vec_63_bits[44], vec_63_bits[29] );
    foobar f1407( dummy[1407], vec_63_bits[45], vec_63_bits[29] );
    foobar f1408( dummy[1408], vec_63_bits[46], vec_63_bits[29] );
    foobar f1409( dummy[1409], vec_63_bits[47], vec_63_bits[29] );
    foobar f1410( dummy[1410], vec_63_bits[48], vec_63_bits[29] );
    foobar f1411( dummy[1411], vec_63_bits[49], vec_63_bits[29] );
    foobar f1412( dummy[1412], vec_63_bits[50], vec_63_bits[29] );
    foobar f1413( dummy[1413], vec_63_bits[51], vec_63_bits[29] );
    foobar f1414( dummy[1414], vec_63_bits[52], vec_63_bits[29] );
    foobar f1415( dummy[1415], vec_63_bits[53], vec_63_bits[29] );
    foobar f1416( dummy[1416], vec_63_bits[54], vec_63_bits[29] );
    foobar f1417( dummy[1417], vec_63_bits[55], vec_63_bits[29] );
    foobar f1418( dummy[1418], vec_63_bits[56], vec_63_bits[29] );
    foobar f1419( dummy[1419], vec_63_bits[57], vec_63_bits[29] );
    foobar f1420( dummy[1420], vec_63_bits[58], vec_63_bits[29] );
    foobar f1421( dummy[1421], vec_63_bits[59], vec_63_bits[29] );
    foobar f1422( dummy[1422], vec_63_bits[60], vec_63_bits[29] );
    foobar f1423( dummy[1423], vec_63_bits[61], vec_63_bits[29] );
    foobar f1424( dummy[1424], vec_63_bits[62], vec_63_bits[29] );
    AN64   an29( o[29], {dummy[1392], dummy[1393], dummy[1394], dummy[1395], dummy[1396], dummy[1397], dummy[1398], dummy[1399], dummy[1400], dummy[1401], dummy[1402], dummy[1403], dummy[1404], dummy[1405], dummy[1406], dummy[1407], dummy[1408], dummy[1409], dummy[1410], dummy[1411], dummy[1412], dummy[1413], dummy[1414], dummy[1415], dummy[1416], dummy[1417], dummy[1418], dummy[1419], dummy[1420], dummy[1421], dummy[1422], dummy[1423], dummy[1424], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1425( dummy[1425], vec_63_bits[31], vec_63_bits[30] );
    foobar f1426( dummy[1426], vec_63_bits[32], vec_63_bits[30] );
    foobar f1427( dummy[1427], vec_63_bits[33], vec_63_bits[30] );
    foobar f1428( dummy[1428], vec_63_bits[34], vec_63_bits[30] );
    foobar f1429( dummy[1429], vec_63_bits[35], vec_63_bits[30] );
    foobar f1430( dummy[1430], vec_63_bits[36], vec_63_bits[30] );
    foobar f1431( dummy[1431], vec_63_bits[37], vec_63_bits[30] );
    foobar f1432( dummy[1432], vec_63_bits[38], vec_63_bits[30] );
    foobar f1433( dummy[1433], vec_63_bits[39], vec_63_bits[30] );
    foobar f1434( dummy[1434], vec_63_bits[40], vec_63_bits[30] );
    foobar f1435( dummy[1435], vec_63_bits[41], vec_63_bits[30] );
    foobar f1436( dummy[1436], vec_63_bits[42], vec_63_bits[30] );
    foobar f1437( dummy[1437], vec_63_bits[43], vec_63_bits[30] );
    foobar f1438( dummy[1438], vec_63_bits[44], vec_63_bits[30] );
    foobar f1439( dummy[1439], vec_63_bits[45], vec_63_bits[30] );
    foobar f1440( dummy[1440], vec_63_bits[46], vec_63_bits[30] );
    foobar f1441( dummy[1441], vec_63_bits[47], vec_63_bits[30] );
    foobar f1442( dummy[1442], vec_63_bits[48], vec_63_bits[30] );
    foobar f1443( dummy[1443], vec_63_bits[49], vec_63_bits[30] );
    foobar f1444( dummy[1444], vec_63_bits[50], vec_63_bits[30] );
    foobar f1445( dummy[1445], vec_63_bits[51], vec_63_bits[30] );
    foobar f1446( dummy[1446], vec_63_bits[52], vec_63_bits[30] );
    foobar f1447( dummy[1447], vec_63_bits[53], vec_63_bits[30] );
    foobar f1448( dummy[1448], vec_63_bits[54], vec_63_bits[30] );
    foobar f1449( dummy[1449], vec_63_bits[55], vec_63_bits[30] );
    foobar f1450( dummy[1450], vec_63_bits[56], vec_63_bits[30] );
    foobar f1451( dummy[1451], vec_63_bits[57], vec_63_bits[30] );
    foobar f1452( dummy[1452], vec_63_bits[58], vec_63_bits[30] );
    foobar f1453( dummy[1453], vec_63_bits[59], vec_63_bits[30] );
    foobar f1454( dummy[1454], vec_63_bits[60], vec_63_bits[30] );
    foobar f1455( dummy[1455], vec_63_bits[61], vec_63_bits[30] );
    foobar f1456( dummy[1456], vec_63_bits[62], vec_63_bits[30] );
    AN64   an30( o[30], {dummy[1425], dummy[1426], dummy[1427], dummy[1428], dummy[1429], dummy[1430], dummy[1431], dummy[1432], dummy[1433], dummy[1434], dummy[1435], dummy[1436], dummy[1437], dummy[1438], dummy[1439], dummy[1440], dummy[1441], dummy[1442], dummy[1443], dummy[1444], dummy[1445], dummy[1446], dummy[1447], dummy[1448], dummy[1449], dummy[1450], dummy[1451], dummy[1452], dummy[1453], dummy[1454], dummy[1455], dummy[1456], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1457( dummy[1457], vec_63_bits[32], vec_63_bits[31] );
    foobar f1458( dummy[1458], vec_63_bits[33], vec_63_bits[31] );
    foobar f1459( dummy[1459], vec_63_bits[34], vec_63_bits[31] );
    foobar f1460( dummy[1460], vec_63_bits[35], vec_63_bits[31] );
    foobar f1461( dummy[1461], vec_63_bits[36], vec_63_bits[31] );
    foobar f1462( dummy[1462], vec_63_bits[37], vec_63_bits[31] );
    foobar f1463( dummy[1463], vec_63_bits[38], vec_63_bits[31] );
    foobar f1464( dummy[1464], vec_63_bits[39], vec_63_bits[31] );
    foobar f1465( dummy[1465], vec_63_bits[40], vec_63_bits[31] );
    foobar f1466( dummy[1466], vec_63_bits[41], vec_63_bits[31] );
    foobar f1467( dummy[1467], vec_63_bits[42], vec_63_bits[31] );
    foobar f1468( dummy[1468], vec_63_bits[43], vec_63_bits[31] );
    foobar f1469( dummy[1469], vec_63_bits[44], vec_63_bits[31] );
    foobar f1470( dummy[1470], vec_63_bits[45], vec_63_bits[31] );
    foobar f1471( dummy[1471], vec_63_bits[46], vec_63_bits[31] );
    foobar f1472( dummy[1472], vec_63_bits[47], vec_63_bits[31] );
    foobar f1473( dummy[1473], vec_63_bits[48], vec_63_bits[31] );
    foobar f1474( dummy[1474], vec_63_bits[49], vec_63_bits[31] );
    foobar f1475( dummy[1475], vec_63_bits[50], vec_63_bits[31] );
    foobar f1476( dummy[1476], vec_63_bits[51], vec_63_bits[31] );
    foobar f1477( dummy[1477], vec_63_bits[52], vec_63_bits[31] );
    foobar f1478( dummy[1478], vec_63_bits[53], vec_63_bits[31] );
    foobar f1479( dummy[1479], vec_63_bits[54], vec_63_bits[31] );
    foobar f1480( dummy[1480], vec_63_bits[55], vec_63_bits[31] );
    foobar f1481( dummy[1481], vec_63_bits[56], vec_63_bits[31] );
    foobar f1482( dummy[1482], vec_63_bits[57], vec_63_bits[31] );
    foobar f1483( dummy[1483], vec_63_bits[58], vec_63_bits[31] );
    foobar f1484( dummy[1484], vec_63_bits[59], vec_63_bits[31] );
    foobar f1485( dummy[1485], vec_63_bits[60], vec_63_bits[31] );
    foobar f1486( dummy[1486], vec_63_bits[61], vec_63_bits[31] );
    foobar f1487( dummy[1487], vec_63_bits[62], vec_63_bits[31] );
    AN64   an31( o[31], {dummy[1457], dummy[1458], dummy[1459], dummy[1460], dummy[1461], dummy[1462], dummy[1463], dummy[1464], dummy[1465], dummy[1466], dummy[1467], dummy[1468], dummy[1469], dummy[1470], dummy[1471], dummy[1472], dummy[1473], dummy[1474], dummy[1475], dummy[1476], dummy[1477], dummy[1478], dummy[1479], dummy[1480], dummy[1481], dummy[1482], dummy[1483], dummy[1484], dummy[1485], dummy[1486], dummy[1487], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1488( dummy[1488], vec_63_bits[33], vec_63_bits[32] );
    foobar f1489( dummy[1489], vec_63_bits[34], vec_63_bits[32] );
    foobar f1490( dummy[1490], vec_63_bits[35], vec_63_bits[32] );
    foobar f1491( dummy[1491], vec_63_bits[36], vec_63_bits[32] );
    foobar f1492( dummy[1492], vec_63_bits[37], vec_63_bits[32] );
    foobar f1493( dummy[1493], vec_63_bits[38], vec_63_bits[32] );
    foobar f1494( dummy[1494], vec_63_bits[39], vec_63_bits[32] );
    foobar f1495( dummy[1495], vec_63_bits[40], vec_63_bits[32] );
    foobar f1496( dummy[1496], vec_63_bits[41], vec_63_bits[32] );
    foobar f1497( dummy[1497], vec_63_bits[42], vec_63_bits[32] );
    foobar f1498( dummy[1498], vec_63_bits[43], vec_63_bits[32] );
    foobar f1499( dummy[1499], vec_63_bits[44], vec_63_bits[32] );
    foobar f1500( dummy[1500], vec_63_bits[45], vec_63_bits[32] );
    foobar f1501( dummy[1501], vec_63_bits[46], vec_63_bits[32] );
    foobar f1502( dummy[1502], vec_63_bits[47], vec_63_bits[32] );
    foobar f1503( dummy[1503], vec_63_bits[48], vec_63_bits[32] );
    foobar f1504( dummy[1504], vec_63_bits[49], vec_63_bits[32] );
    foobar f1505( dummy[1505], vec_63_bits[50], vec_63_bits[32] );
    foobar f1506( dummy[1506], vec_63_bits[51], vec_63_bits[32] );
    foobar f1507( dummy[1507], vec_63_bits[52], vec_63_bits[32] );
    foobar f1508( dummy[1508], vec_63_bits[53], vec_63_bits[32] );
    foobar f1509( dummy[1509], vec_63_bits[54], vec_63_bits[32] );
    foobar f1510( dummy[1510], vec_63_bits[55], vec_63_bits[32] );
    foobar f1511( dummy[1511], vec_63_bits[56], vec_63_bits[32] );
    foobar f1512( dummy[1512], vec_63_bits[57], vec_63_bits[32] );
    foobar f1513( dummy[1513], vec_63_bits[58], vec_63_bits[32] );
    foobar f1514( dummy[1514], vec_63_bits[59], vec_63_bits[32] );
    foobar f1515( dummy[1515], vec_63_bits[60], vec_63_bits[32] );
    foobar f1516( dummy[1516], vec_63_bits[61], vec_63_bits[32] );
    foobar f1517( dummy[1517], vec_63_bits[62], vec_63_bits[32] );
    AN64   an32( o[32], {dummy[1488], dummy[1489], dummy[1490], dummy[1491], dummy[1492], dummy[1493], dummy[1494], dummy[1495], dummy[1496], dummy[1497], dummy[1498], dummy[1499], dummy[1500], dummy[1501], dummy[1502], dummy[1503], dummy[1504], dummy[1505], dummy[1506], dummy[1507], dummy[1508], dummy[1509], dummy[1510], dummy[1511], dummy[1512], dummy[1513], dummy[1514], dummy[1515], dummy[1516], dummy[1517], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1518( dummy[1518], vec_63_bits[34], vec_63_bits[33] );
    foobar f1519( dummy[1519], vec_63_bits[35], vec_63_bits[33] );
    foobar f1520( dummy[1520], vec_63_bits[36], vec_63_bits[33] );
    foobar f1521( dummy[1521], vec_63_bits[37], vec_63_bits[33] );
    foobar f1522( dummy[1522], vec_63_bits[38], vec_63_bits[33] );
    foobar f1523( dummy[1523], vec_63_bits[39], vec_63_bits[33] );
    foobar f1524( dummy[1524], vec_63_bits[40], vec_63_bits[33] );
    foobar f1525( dummy[1525], vec_63_bits[41], vec_63_bits[33] );
    foobar f1526( dummy[1526], vec_63_bits[42], vec_63_bits[33] );
    foobar f1527( dummy[1527], vec_63_bits[43], vec_63_bits[33] );
    foobar f1528( dummy[1528], vec_63_bits[44], vec_63_bits[33] );
    foobar f1529( dummy[1529], vec_63_bits[45], vec_63_bits[33] );
    foobar f1530( dummy[1530], vec_63_bits[46], vec_63_bits[33] );
    foobar f1531( dummy[1531], vec_63_bits[47], vec_63_bits[33] );
    foobar f1532( dummy[1532], vec_63_bits[48], vec_63_bits[33] );
    foobar f1533( dummy[1533], vec_63_bits[49], vec_63_bits[33] );
    foobar f1534( dummy[1534], vec_63_bits[50], vec_63_bits[33] );
    foobar f1535( dummy[1535], vec_63_bits[51], vec_63_bits[33] );
    foobar f1536( dummy[1536], vec_63_bits[52], vec_63_bits[33] );
    foobar f1537( dummy[1537], vec_63_bits[53], vec_63_bits[33] );
    foobar f1538( dummy[1538], vec_63_bits[54], vec_63_bits[33] );
    foobar f1539( dummy[1539], vec_63_bits[55], vec_63_bits[33] );
    foobar f1540( dummy[1540], vec_63_bits[56], vec_63_bits[33] );
    foobar f1541( dummy[1541], vec_63_bits[57], vec_63_bits[33] );
    foobar f1542( dummy[1542], vec_63_bits[58], vec_63_bits[33] );
    foobar f1543( dummy[1543], vec_63_bits[59], vec_63_bits[33] );
    foobar f1544( dummy[1544], vec_63_bits[60], vec_63_bits[33] );
    foobar f1545( dummy[1545], vec_63_bits[61], vec_63_bits[33] );
    foobar f1546( dummy[1546], vec_63_bits[62], vec_63_bits[33] );
    AN64   an33( o[33], {dummy[1518], dummy[1519], dummy[1520], dummy[1521], dummy[1522], dummy[1523], dummy[1524], dummy[1525], dummy[1526], dummy[1527], dummy[1528], dummy[1529], dummy[1530], dummy[1531], dummy[1532], dummy[1533], dummy[1534], dummy[1535], dummy[1536], dummy[1537], dummy[1538], dummy[1539], dummy[1540], dummy[1541], dummy[1542], dummy[1543], dummy[1544], dummy[1545], dummy[1546], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1547( dummy[1547], vec_63_bits[35], vec_63_bits[34] );
    foobar f1548( dummy[1548], vec_63_bits[36], vec_63_bits[34] );
    foobar f1549( dummy[1549], vec_63_bits[37], vec_63_bits[34] );
    foobar f1550( dummy[1550], vec_63_bits[38], vec_63_bits[34] );
    foobar f1551( dummy[1551], vec_63_bits[39], vec_63_bits[34] );
    foobar f1552( dummy[1552], vec_63_bits[40], vec_63_bits[34] );
    foobar f1553( dummy[1553], vec_63_bits[41], vec_63_bits[34] );
    foobar f1554( dummy[1554], vec_63_bits[42], vec_63_bits[34] );
    foobar f1555( dummy[1555], vec_63_bits[43], vec_63_bits[34] );
    foobar f1556( dummy[1556], vec_63_bits[44], vec_63_bits[34] );
    foobar f1557( dummy[1557], vec_63_bits[45], vec_63_bits[34] );
    foobar f1558( dummy[1558], vec_63_bits[46], vec_63_bits[34] );
    foobar f1559( dummy[1559], vec_63_bits[47], vec_63_bits[34] );
    foobar f1560( dummy[1560], vec_63_bits[48], vec_63_bits[34] );
    foobar f1561( dummy[1561], vec_63_bits[49], vec_63_bits[34] );
    foobar f1562( dummy[1562], vec_63_bits[50], vec_63_bits[34] );
    foobar f1563( dummy[1563], vec_63_bits[51], vec_63_bits[34] );
    foobar f1564( dummy[1564], vec_63_bits[52], vec_63_bits[34] );
    foobar f1565( dummy[1565], vec_63_bits[53], vec_63_bits[34] );
    foobar f1566( dummy[1566], vec_63_bits[54], vec_63_bits[34] );
    foobar f1567( dummy[1567], vec_63_bits[55], vec_63_bits[34] );
    foobar f1568( dummy[1568], vec_63_bits[56], vec_63_bits[34] );
    foobar f1569( dummy[1569], vec_63_bits[57], vec_63_bits[34] );
    foobar f1570( dummy[1570], vec_63_bits[58], vec_63_bits[34] );
    foobar f1571( dummy[1571], vec_63_bits[59], vec_63_bits[34] );
    foobar f1572( dummy[1572], vec_63_bits[60], vec_63_bits[34] );
    foobar f1573( dummy[1573], vec_63_bits[61], vec_63_bits[34] );
    foobar f1574( dummy[1574], vec_63_bits[62], vec_63_bits[34] );
    AN64   an34( o[34], {dummy[1547], dummy[1548], dummy[1549], dummy[1550], dummy[1551], dummy[1552], dummy[1553], dummy[1554], dummy[1555], dummy[1556], dummy[1557], dummy[1558], dummy[1559], dummy[1560], dummy[1561], dummy[1562], dummy[1563], dummy[1564], dummy[1565], dummy[1566], dummy[1567], dummy[1568], dummy[1569], dummy[1570], dummy[1571], dummy[1572], dummy[1573], dummy[1574], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1575( dummy[1575], vec_63_bits[36], vec_63_bits[35] );
    foobar f1576( dummy[1576], vec_63_bits[37], vec_63_bits[35] );
    foobar f1577( dummy[1577], vec_63_bits[38], vec_63_bits[35] );
    foobar f1578( dummy[1578], vec_63_bits[39], vec_63_bits[35] );
    foobar f1579( dummy[1579], vec_63_bits[40], vec_63_bits[35] );
    foobar f1580( dummy[1580], vec_63_bits[41], vec_63_bits[35] );
    foobar f1581( dummy[1581], vec_63_bits[42], vec_63_bits[35] );
    foobar f1582( dummy[1582], vec_63_bits[43], vec_63_bits[35] );
    foobar f1583( dummy[1583], vec_63_bits[44], vec_63_bits[35] );
    foobar f1584( dummy[1584], vec_63_bits[45], vec_63_bits[35] );
    foobar f1585( dummy[1585], vec_63_bits[46], vec_63_bits[35] );
    foobar f1586( dummy[1586], vec_63_bits[47], vec_63_bits[35] );
    foobar f1587( dummy[1587], vec_63_bits[48], vec_63_bits[35] );
    foobar f1588( dummy[1588], vec_63_bits[49], vec_63_bits[35] );
    foobar f1589( dummy[1589], vec_63_bits[50], vec_63_bits[35] );
    foobar f1590( dummy[1590], vec_63_bits[51], vec_63_bits[35] );
    foobar f1591( dummy[1591], vec_63_bits[52], vec_63_bits[35] );
    foobar f1592( dummy[1592], vec_63_bits[53], vec_63_bits[35] );
    foobar f1593( dummy[1593], vec_63_bits[54], vec_63_bits[35] );
    foobar f1594( dummy[1594], vec_63_bits[55], vec_63_bits[35] );
    foobar f1595( dummy[1595], vec_63_bits[56], vec_63_bits[35] );
    foobar f1596( dummy[1596], vec_63_bits[57], vec_63_bits[35] );
    foobar f1597( dummy[1597], vec_63_bits[58], vec_63_bits[35] );
    foobar f1598( dummy[1598], vec_63_bits[59], vec_63_bits[35] );
    foobar f1599( dummy[1599], vec_63_bits[60], vec_63_bits[35] );
    foobar f1600( dummy[1600], vec_63_bits[61], vec_63_bits[35] );
    foobar f1601( dummy[1601], vec_63_bits[62], vec_63_bits[35] );
    AN64   an35( o[35], {dummy[1575], dummy[1576], dummy[1577], dummy[1578], dummy[1579], dummy[1580], dummy[1581], dummy[1582], dummy[1583], dummy[1584], dummy[1585], dummy[1586], dummy[1587], dummy[1588], dummy[1589], dummy[1590], dummy[1591], dummy[1592], dummy[1593], dummy[1594], dummy[1595], dummy[1596], dummy[1597], dummy[1598], dummy[1599], dummy[1600], dummy[1601], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1602( dummy[1602], vec_63_bits[37], vec_63_bits[36] );
    foobar f1603( dummy[1603], vec_63_bits[38], vec_63_bits[36] );
    foobar f1604( dummy[1604], vec_63_bits[39], vec_63_bits[36] );
    foobar f1605( dummy[1605], vec_63_bits[40], vec_63_bits[36] );
    foobar f1606( dummy[1606], vec_63_bits[41], vec_63_bits[36] );
    foobar f1607( dummy[1607], vec_63_bits[42], vec_63_bits[36] );
    foobar f1608( dummy[1608], vec_63_bits[43], vec_63_bits[36] );
    foobar f1609( dummy[1609], vec_63_bits[44], vec_63_bits[36] );
    foobar f1610( dummy[1610], vec_63_bits[45], vec_63_bits[36] );
    foobar f1611( dummy[1611], vec_63_bits[46], vec_63_bits[36] );
    foobar f1612( dummy[1612], vec_63_bits[47], vec_63_bits[36] );
    foobar f1613( dummy[1613], vec_63_bits[48], vec_63_bits[36] );
    foobar f1614( dummy[1614], vec_63_bits[49], vec_63_bits[36] );
    foobar f1615( dummy[1615], vec_63_bits[50], vec_63_bits[36] );
    foobar f1616( dummy[1616], vec_63_bits[51], vec_63_bits[36] );
    foobar f1617( dummy[1617], vec_63_bits[52], vec_63_bits[36] );
    foobar f1618( dummy[1618], vec_63_bits[53], vec_63_bits[36] );
    foobar f1619( dummy[1619], vec_63_bits[54], vec_63_bits[36] );
    foobar f1620( dummy[1620], vec_63_bits[55], vec_63_bits[36] );
    foobar f1621( dummy[1621], vec_63_bits[56], vec_63_bits[36] );
    foobar f1622( dummy[1622], vec_63_bits[57], vec_63_bits[36] );
    foobar f1623( dummy[1623], vec_63_bits[58], vec_63_bits[36] );
    foobar f1624( dummy[1624], vec_63_bits[59], vec_63_bits[36] );
    foobar f1625( dummy[1625], vec_63_bits[60], vec_63_bits[36] );
    foobar f1626( dummy[1626], vec_63_bits[61], vec_63_bits[36] );
    foobar f1627( dummy[1627], vec_63_bits[62], vec_63_bits[36] );
    AN64   an36( o[36], {dummy[1602], dummy[1603], dummy[1604], dummy[1605], dummy[1606], dummy[1607], dummy[1608], dummy[1609], dummy[1610], dummy[1611], dummy[1612], dummy[1613], dummy[1614], dummy[1615], dummy[1616], dummy[1617], dummy[1618], dummy[1619], dummy[1620], dummy[1621], dummy[1622], dummy[1623], dummy[1624], dummy[1625], dummy[1626], dummy[1627], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1628( dummy[1628], vec_63_bits[38], vec_63_bits[37] );
    foobar f1629( dummy[1629], vec_63_bits[39], vec_63_bits[37] );
    foobar f1630( dummy[1630], vec_63_bits[40], vec_63_bits[37] );
    foobar f1631( dummy[1631], vec_63_bits[41], vec_63_bits[37] );
    foobar f1632( dummy[1632], vec_63_bits[42], vec_63_bits[37] );
    foobar f1633( dummy[1633], vec_63_bits[43], vec_63_bits[37] );
    foobar f1634( dummy[1634], vec_63_bits[44], vec_63_bits[37] );
    foobar f1635( dummy[1635], vec_63_bits[45], vec_63_bits[37] );
    foobar f1636( dummy[1636], vec_63_bits[46], vec_63_bits[37] );
    foobar f1637( dummy[1637], vec_63_bits[47], vec_63_bits[37] );
    foobar f1638( dummy[1638], vec_63_bits[48], vec_63_bits[37] );
    foobar f1639( dummy[1639], vec_63_bits[49], vec_63_bits[37] );
    foobar f1640( dummy[1640], vec_63_bits[50], vec_63_bits[37] );
    foobar f1641( dummy[1641], vec_63_bits[51], vec_63_bits[37] );
    foobar f1642( dummy[1642], vec_63_bits[52], vec_63_bits[37] );
    foobar f1643( dummy[1643], vec_63_bits[53], vec_63_bits[37] );
    foobar f1644( dummy[1644], vec_63_bits[54], vec_63_bits[37] );
    foobar f1645( dummy[1645], vec_63_bits[55], vec_63_bits[37] );
    foobar f1646( dummy[1646], vec_63_bits[56], vec_63_bits[37] );
    foobar f1647( dummy[1647], vec_63_bits[57], vec_63_bits[37] );
    foobar f1648( dummy[1648], vec_63_bits[58], vec_63_bits[37] );
    foobar f1649( dummy[1649], vec_63_bits[59], vec_63_bits[37] );
    foobar f1650( dummy[1650], vec_63_bits[60], vec_63_bits[37] );
    foobar f1651( dummy[1651], vec_63_bits[61], vec_63_bits[37] );
    foobar f1652( dummy[1652], vec_63_bits[62], vec_63_bits[37] );
    AN64   an37( o[37], {dummy[1628], dummy[1629], dummy[1630], dummy[1631], dummy[1632], dummy[1633], dummy[1634], dummy[1635], dummy[1636], dummy[1637], dummy[1638], dummy[1639], dummy[1640], dummy[1641], dummy[1642], dummy[1643], dummy[1644], dummy[1645], dummy[1646], dummy[1647], dummy[1648], dummy[1649], dummy[1650], dummy[1651], dummy[1652], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1653( dummy[1653], vec_63_bits[39], vec_63_bits[38] );
    foobar f1654( dummy[1654], vec_63_bits[40], vec_63_bits[38] );
    foobar f1655( dummy[1655], vec_63_bits[41], vec_63_bits[38] );
    foobar f1656( dummy[1656], vec_63_bits[42], vec_63_bits[38] );
    foobar f1657( dummy[1657], vec_63_bits[43], vec_63_bits[38] );
    foobar f1658( dummy[1658], vec_63_bits[44], vec_63_bits[38] );
    foobar f1659( dummy[1659], vec_63_bits[45], vec_63_bits[38] );
    foobar f1660( dummy[1660], vec_63_bits[46], vec_63_bits[38] );
    foobar f1661( dummy[1661], vec_63_bits[47], vec_63_bits[38] );
    foobar f1662( dummy[1662], vec_63_bits[48], vec_63_bits[38] );
    foobar f1663( dummy[1663], vec_63_bits[49], vec_63_bits[38] );
    foobar f1664( dummy[1664], vec_63_bits[50], vec_63_bits[38] );
    foobar f1665( dummy[1665], vec_63_bits[51], vec_63_bits[38] );
    foobar f1666( dummy[1666], vec_63_bits[52], vec_63_bits[38] );
    foobar f1667( dummy[1667], vec_63_bits[53], vec_63_bits[38] );
    foobar f1668( dummy[1668], vec_63_bits[54], vec_63_bits[38] );
    foobar f1669( dummy[1669], vec_63_bits[55], vec_63_bits[38] );
    foobar f1670( dummy[1670], vec_63_bits[56], vec_63_bits[38] );
    foobar f1671( dummy[1671], vec_63_bits[57], vec_63_bits[38] );
    foobar f1672( dummy[1672], vec_63_bits[58], vec_63_bits[38] );
    foobar f1673( dummy[1673], vec_63_bits[59], vec_63_bits[38] );
    foobar f1674( dummy[1674], vec_63_bits[60], vec_63_bits[38] );
    foobar f1675( dummy[1675], vec_63_bits[61], vec_63_bits[38] );
    foobar f1676( dummy[1676], vec_63_bits[62], vec_63_bits[38] );
    AN64   an38( o[38], {dummy[1653], dummy[1654], dummy[1655], dummy[1656], dummy[1657], dummy[1658], dummy[1659], dummy[1660], dummy[1661], dummy[1662], dummy[1663], dummy[1664], dummy[1665], dummy[1666], dummy[1667], dummy[1668], dummy[1669], dummy[1670], dummy[1671], dummy[1672], dummy[1673], dummy[1674], dummy[1675], dummy[1676], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1677( dummy[1677], vec_63_bits[40], vec_63_bits[39] );
    foobar f1678( dummy[1678], vec_63_bits[41], vec_63_bits[39] );
    foobar f1679( dummy[1679], vec_63_bits[42], vec_63_bits[39] );
    foobar f1680( dummy[1680], vec_63_bits[43], vec_63_bits[39] );
    foobar f1681( dummy[1681], vec_63_bits[44], vec_63_bits[39] );
    foobar f1682( dummy[1682], vec_63_bits[45], vec_63_bits[39] );
    foobar f1683( dummy[1683], vec_63_bits[46], vec_63_bits[39] );
    foobar f1684( dummy[1684], vec_63_bits[47], vec_63_bits[39] );
    foobar f1685( dummy[1685], vec_63_bits[48], vec_63_bits[39] );
    foobar f1686( dummy[1686], vec_63_bits[49], vec_63_bits[39] );
    foobar f1687( dummy[1687], vec_63_bits[50], vec_63_bits[39] );
    foobar f1688( dummy[1688], vec_63_bits[51], vec_63_bits[39] );
    foobar f1689( dummy[1689], vec_63_bits[52], vec_63_bits[39] );
    foobar f1690( dummy[1690], vec_63_bits[53], vec_63_bits[39] );
    foobar f1691( dummy[1691], vec_63_bits[54], vec_63_bits[39] );
    foobar f1692( dummy[1692], vec_63_bits[55], vec_63_bits[39] );
    foobar f1693( dummy[1693], vec_63_bits[56], vec_63_bits[39] );
    foobar f1694( dummy[1694], vec_63_bits[57], vec_63_bits[39] );
    foobar f1695( dummy[1695], vec_63_bits[58], vec_63_bits[39] );
    foobar f1696( dummy[1696], vec_63_bits[59], vec_63_bits[39] );
    foobar f1697( dummy[1697], vec_63_bits[60], vec_63_bits[39] );
    foobar f1698( dummy[1698], vec_63_bits[61], vec_63_bits[39] );
    foobar f1699( dummy[1699], vec_63_bits[62], vec_63_bits[39] );
    AN64   an39( o[39], {dummy[1677], dummy[1678], dummy[1679], dummy[1680], dummy[1681], dummy[1682], dummy[1683], dummy[1684], dummy[1685], dummy[1686], dummy[1687], dummy[1688], dummy[1689], dummy[1690], dummy[1691], dummy[1692], dummy[1693], dummy[1694], dummy[1695], dummy[1696], dummy[1697], dummy[1698], dummy[1699], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1700( dummy[1700], vec_63_bits[41], vec_63_bits[40] );
    foobar f1701( dummy[1701], vec_63_bits[42], vec_63_bits[40] );
    foobar f1702( dummy[1702], vec_63_bits[43], vec_63_bits[40] );
    foobar f1703( dummy[1703], vec_63_bits[44], vec_63_bits[40] );
    foobar f1704( dummy[1704], vec_63_bits[45], vec_63_bits[40] );
    foobar f1705( dummy[1705], vec_63_bits[46], vec_63_bits[40] );
    foobar f1706( dummy[1706], vec_63_bits[47], vec_63_bits[40] );
    foobar f1707( dummy[1707], vec_63_bits[48], vec_63_bits[40] );
    foobar f1708( dummy[1708], vec_63_bits[49], vec_63_bits[40] );
    foobar f1709( dummy[1709], vec_63_bits[50], vec_63_bits[40] );
    foobar f1710( dummy[1710], vec_63_bits[51], vec_63_bits[40] );
    foobar f1711( dummy[1711], vec_63_bits[52], vec_63_bits[40] );
    foobar f1712( dummy[1712], vec_63_bits[53], vec_63_bits[40] );
    foobar f1713( dummy[1713], vec_63_bits[54], vec_63_bits[40] );
    foobar f1714( dummy[1714], vec_63_bits[55], vec_63_bits[40] );
    foobar f1715( dummy[1715], vec_63_bits[56], vec_63_bits[40] );
    foobar f1716( dummy[1716], vec_63_bits[57], vec_63_bits[40] );
    foobar f1717( dummy[1717], vec_63_bits[58], vec_63_bits[40] );
    foobar f1718( dummy[1718], vec_63_bits[59], vec_63_bits[40] );
    foobar f1719( dummy[1719], vec_63_bits[60], vec_63_bits[40] );
    foobar f1720( dummy[1720], vec_63_bits[61], vec_63_bits[40] );
    foobar f1721( dummy[1721], vec_63_bits[62], vec_63_bits[40] );
    AN64   an40( o[40], {dummy[1700], dummy[1701], dummy[1702], dummy[1703], dummy[1704], dummy[1705], dummy[1706], dummy[1707], dummy[1708], dummy[1709], dummy[1710], dummy[1711], dummy[1712], dummy[1713], dummy[1714], dummy[1715], dummy[1716], dummy[1717], dummy[1718], dummy[1719], dummy[1720], dummy[1721], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1722( dummy[1722], vec_63_bits[42], vec_63_bits[41] );
    foobar f1723( dummy[1723], vec_63_bits[43], vec_63_bits[41] );
    foobar f1724( dummy[1724], vec_63_bits[44], vec_63_bits[41] );
    foobar f1725( dummy[1725], vec_63_bits[45], vec_63_bits[41] );
    foobar f1726( dummy[1726], vec_63_bits[46], vec_63_bits[41] );
    foobar f1727( dummy[1727], vec_63_bits[47], vec_63_bits[41] );
    foobar f1728( dummy[1728], vec_63_bits[48], vec_63_bits[41] );
    foobar f1729( dummy[1729], vec_63_bits[49], vec_63_bits[41] );
    foobar f1730( dummy[1730], vec_63_bits[50], vec_63_bits[41] );
    foobar f1731( dummy[1731], vec_63_bits[51], vec_63_bits[41] );
    foobar f1732( dummy[1732], vec_63_bits[52], vec_63_bits[41] );
    foobar f1733( dummy[1733], vec_63_bits[53], vec_63_bits[41] );
    foobar f1734( dummy[1734], vec_63_bits[54], vec_63_bits[41] );
    foobar f1735( dummy[1735], vec_63_bits[55], vec_63_bits[41] );
    foobar f1736( dummy[1736], vec_63_bits[56], vec_63_bits[41] );
    foobar f1737( dummy[1737], vec_63_bits[57], vec_63_bits[41] );
    foobar f1738( dummy[1738], vec_63_bits[58], vec_63_bits[41] );
    foobar f1739( dummy[1739], vec_63_bits[59], vec_63_bits[41] );
    foobar f1740( dummy[1740], vec_63_bits[60], vec_63_bits[41] );
    foobar f1741( dummy[1741], vec_63_bits[61], vec_63_bits[41] );
    foobar f1742( dummy[1742], vec_63_bits[62], vec_63_bits[41] );
    AN64   an41( o[41], {dummy[1722], dummy[1723], dummy[1724], dummy[1725], dummy[1726], dummy[1727], dummy[1728], dummy[1729], dummy[1730], dummy[1731], dummy[1732], dummy[1733], dummy[1734], dummy[1735], dummy[1736], dummy[1737], dummy[1738], dummy[1739], dummy[1740], dummy[1741], dummy[1742], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1743( dummy[1743], vec_63_bits[43], vec_63_bits[42] );
    foobar f1744( dummy[1744], vec_63_bits[44], vec_63_bits[42] );
    foobar f1745( dummy[1745], vec_63_bits[45], vec_63_bits[42] );
    foobar f1746( dummy[1746], vec_63_bits[46], vec_63_bits[42] );
    foobar f1747( dummy[1747], vec_63_bits[47], vec_63_bits[42] );
    foobar f1748( dummy[1748], vec_63_bits[48], vec_63_bits[42] );
    foobar f1749( dummy[1749], vec_63_bits[49], vec_63_bits[42] );
    foobar f1750( dummy[1750], vec_63_bits[50], vec_63_bits[42] );
    foobar f1751( dummy[1751], vec_63_bits[51], vec_63_bits[42] );
    foobar f1752( dummy[1752], vec_63_bits[52], vec_63_bits[42] );
    foobar f1753( dummy[1753], vec_63_bits[53], vec_63_bits[42] );
    foobar f1754( dummy[1754], vec_63_bits[54], vec_63_bits[42] );
    foobar f1755( dummy[1755], vec_63_bits[55], vec_63_bits[42] );
    foobar f1756( dummy[1756], vec_63_bits[56], vec_63_bits[42] );
    foobar f1757( dummy[1757], vec_63_bits[57], vec_63_bits[42] );
    foobar f1758( dummy[1758], vec_63_bits[58], vec_63_bits[42] );
    foobar f1759( dummy[1759], vec_63_bits[59], vec_63_bits[42] );
    foobar f1760( dummy[1760], vec_63_bits[60], vec_63_bits[42] );
    foobar f1761( dummy[1761], vec_63_bits[61], vec_63_bits[42] );
    foobar f1762( dummy[1762], vec_63_bits[62], vec_63_bits[42] );
    AN64   an42( o[42], {dummy[1743], dummy[1744], dummy[1745], dummy[1746], dummy[1747], dummy[1748], dummy[1749], dummy[1750], dummy[1751], dummy[1752], dummy[1753], dummy[1754], dummy[1755], dummy[1756], dummy[1757], dummy[1758], dummy[1759], dummy[1760], dummy[1761], dummy[1762], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1763( dummy[1763], vec_63_bits[44], vec_63_bits[43] );
    foobar f1764( dummy[1764], vec_63_bits[45], vec_63_bits[43] );
    foobar f1765( dummy[1765], vec_63_bits[46], vec_63_bits[43] );
    foobar f1766( dummy[1766], vec_63_bits[47], vec_63_bits[43] );
    foobar f1767( dummy[1767], vec_63_bits[48], vec_63_bits[43] );
    foobar f1768( dummy[1768], vec_63_bits[49], vec_63_bits[43] );
    foobar f1769( dummy[1769], vec_63_bits[50], vec_63_bits[43] );
    foobar f1770( dummy[1770], vec_63_bits[51], vec_63_bits[43] );
    foobar f1771( dummy[1771], vec_63_bits[52], vec_63_bits[43] );
    foobar f1772( dummy[1772], vec_63_bits[53], vec_63_bits[43] );
    foobar f1773( dummy[1773], vec_63_bits[54], vec_63_bits[43] );
    foobar f1774( dummy[1774], vec_63_bits[55], vec_63_bits[43] );
    foobar f1775( dummy[1775], vec_63_bits[56], vec_63_bits[43] );
    foobar f1776( dummy[1776], vec_63_bits[57], vec_63_bits[43] );
    foobar f1777( dummy[1777], vec_63_bits[58], vec_63_bits[43] );
    foobar f1778( dummy[1778], vec_63_bits[59], vec_63_bits[43] );
    foobar f1779( dummy[1779], vec_63_bits[60], vec_63_bits[43] );
    foobar f1780( dummy[1780], vec_63_bits[61], vec_63_bits[43] );
    foobar f1781( dummy[1781], vec_63_bits[62], vec_63_bits[43] );
    AN64   an43( o[43], {dummy[1763], dummy[1764], dummy[1765], dummy[1766], dummy[1767], dummy[1768], dummy[1769], dummy[1770], dummy[1771], dummy[1772], dummy[1773], dummy[1774], dummy[1775], dummy[1776], dummy[1777], dummy[1778], dummy[1779], dummy[1780], dummy[1781], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1782( dummy[1782], vec_63_bits[45], vec_63_bits[44] );
    foobar f1783( dummy[1783], vec_63_bits[46], vec_63_bits[44] );
    foobar f1784( dummy[1784], vec_63_bits[47], vec_63_bits[44] );
    foobar f1785( dummy[1785], vec_63_bits[48], vec_63_bits[44] );
    foobar f1786( dummy[1786], vec_63_bits[49], vec_63_bits[44] );
    foobar f1787( dummy[1787], vec_63_bits[50], vec_63_bits[44] );
    foobar f1788( dummy[1788], vec_63_bits[51], vec_63_bits[44] );
    foobar f1789( dummy[1789], vec_63_bits[52], vec_63_bits[44] );
    foobar f1790( dummy[1790], vec_63_bits[53], vec_63_bits[44] );
    foobar f1791( dummy[1791], vec_63_bits[54], vec_63_bits[44] );
    foobar f1792( dummy[1792], vec_63_bits[55], vec_63_bits[44] );
    foobar f1793( dummy[1793], vec_63_bits[56], vec_63_bits[44] );
    foobar f1794( dummy[1794], vec_63_bits[57], vec_63_bits[44] );
    foobar f1795( dummy[1795], vec_63_bits[58], vec_63_bits[44] );
    foobar f1796( dummy[1796], vec_63_bits[59], vec_63_bits[44] );
    foobar f1797( dummy[1797], vec_63_bits[60], vec_63_bits[44] );
    foobar f1798( dummy[1798], vec_63_bits[61], vec_63_bits[44] );
    foobar f1799( dummy[1799], vec_63_bits[62], vec_63_bits[44] );
    AN64   an44( o[44], {dummy[1782], dummy[1783], dummy[1784], dummy[1785], dummy[1786], dummy[1787], dummy[1788], dummy[1789], dummy[1790], dummy[1791], dummy[1792], dummy[1793], dummy[1794], dummy[1795], dummy[1796], dummy[1797], dummy[1798], dummy[1799], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1800( dummy[1800], vec_63_bits[46], vec_63_bits[45] );
    foobar f1801( dummy[1801], vec_63_bits[47], vec_63_bits[45] );
    foobar f1802( dummy[1802], vec_63_bits[48], vec_63_bits[45] );
    foobar f1803( dummy[1803], vec_63_bits[49], vec_63_bits[45] );
    foobar f1804( dummy[1804], vec_63_bits[50], vec_63_bits[45] );
    foobar f1805( dummy[1805], vec_63_bits[51], vec_63_bits[45] );
    foobar f1806( dummy[1806], vec_63_bits[52], vec_63_bits[45] );
    foobar f1807( dummy[1807], vec_63_bits[53], vec_63_bits[45] );
    foobar f1808( dummy[1808], vec_63_bits[54], vec_63_bits[45] );
    foobar f1809( dummy[1809], vec_63_bits[55], vec_63_bits[45] );
    foobar f1810( dummy[1810], vec_63_bits[56], vec_63_bits[45] );
    foobar f1811( dummy[1811], vec_63_bits[57], vec_63_bits[45] );
    foobar f1812( dummy[1812], vec_63_bits[58], vec_63_bits[45] );
    foobar f1813( dummy[1813], vec_63_bits[59], vec_63_bits[45] );
    foobar f1814( dummy[1814], vec_63_bits[60], vec_63_bits[45] );
    foobar f1815( dummy[1815], vec_63_bits[61], vec_63_bits[45] );
    foobar f1816( dummy[1816], vec_63_bits[62], vec_63_bits[45] );
    AN64   an45( o[45], {dummy[1800], dummy[1801], dummy[1802], dummy[1803], dummy[1804], dummy[1805], dummy[1806], dummy[1807], dummy[1808], dummy[1809], dummy[1810], dummy[1811], dummy[1812], dummy[1813], dummy[1814], dummy[1815], dummy[1816], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1817( dummy[1817], vec_63_bits[47], vec_63_bits[46] );
    foobar f1818( dummy[1818], vec_63_bits[48], vec_63_bits[46] );
    foobar f1819( dummy[1819], vec_63_bits[49], vec_63_bits[46] );
    foobar f1820( dummy[1820], vec_63_bits[50], vec_63_bits[46] );
    foobar f1821( dummy[1821], vec_63_bits[51], vec_63_bits[46] );
    foobar f1822( dummy[1822], vec_63_bits[52], vec_63_bits[46] );
    foobar f1823( dummy[1823], vec_63_bits[53], vec_63_bits[46] );
    foobar f1824( dummy[1824], vec_63_bits[54], vec_63_bits[46] );
    foobar f1825( dummy[1825], vec_63_bits[55], vec_63_bits[46] );
    foobar f1826( dummy[1826], vec_63_bits[56], vec_63_bits[46] );
    foobar f1827( dummy[1827], vec_63_bits[57], vec_63_bits[46] );
    foobar f1828( dummy[1828], vec_63_bits[58], vec_63_bits[46] );
    foobar f1829( dummy[1829], vec_63_bits[59], vec_63_bits[46] );
    foobar f1830( dummy[1830], vec_63_bits[60], vec_63_bits[46] );
    foobar f1831( dummy[1831], vec_63_bits[61], vec_63_bits[46] );
    foobar f1832( dummy[1832], vec_63_bits[62], vec_63_bits[46] );
    AN64   an46( o[46], {dummy[1817], dummy[1818], dummy[1819], dummy[1820], dummy[1821], dummy[1822], dummy[1823], dummy[1824], dummy[1825], dummy[1826], dummy[1827], dummy[1828], dummy[1829], dummy[1830], dummy[1831], dummy[1832], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1833( dummy[1833], vec_63_bits[48], vec_63_bits[47] );
    foobar f1834( dummy[1834], vec_63_bits[49], vec_63_bits[47] );
    foobar f1835( dummy[1835], vec_63_bits[50], vec_63_bits[47] );
    foobar f1836( dummy[1836], vec_63_bits[51], vec_63_bits[47] );
    foobar f1837( dummy[1837], vec_63_bits[52], vec_63_bits[47] );
    foobar f1838( dummy[1838], vec_63_bits[53], vec_63_bits[47] );
    foobar f1839( dummy[1839], vec_63_bits[54], vec_63_bits[47] );
    foobar f1840( dummy[1840], vec_63_bits[55], vec_63_bits[47] );
    foobar f1841( dummy[1841], vec_63_bits[56], vec_63_bits[47] );
    foobar f1842( dummy[1842], vec_63_bits[57], vec_63_bits[47] );
    foobar f1843( dummy[1843], vec_63_bits[58], vec_63_bits[47] );
    foobar f1844( dummy[1844], vec_63_bits[59], vec_63_bits[47] );
    foobar f1845( dummy[1845], vec_63_bits[60], vec_63_bits[47] );
    foobar f1846( dummy[1846], vec_63_bits[61], vec_63_bits[47] );
    foobar f1847( dummy[1847], vec_63_bits[62], vec_63_bits[47] );
    AN64   an47( o[47], {dummy[1833], dummy[1834], dummy[1835], dummy[1836], dummy[1837], dummy[1838], dummy[1839], dummy[1840], dummy[1841], dummy[1842], dummy[1843], dummy[1844], dummy[1845], dummy[1846], dummy[1847], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1848( dummy[1848], vec_63_bits[49], vec_63_bits[48] );
    foobar f1849( dummy[1849], vec_63_bits[50], vec_63_bits[48] );
    foobar f1850( dummy[1850], vec_63_bits[51], vec_63_bits[48] );
    foobar f1851( dummy[1851], vec_63_bits[52], vec_63_bits[48] );
    foobar f1852( dummy[1852], vec_63_bits[53], vec_63_bits[48] );
    foobar f1853( dummy[1853], vec_63_bits[54], vec_63_bits[48] );
    foobar f1854( dummy[1854], vec_63_bits[55], vec_63_bits[48] );
    foobar f1855( dummy[1855], vec_63_bits[56], vec_63_bits[48] );
    foobar f1856( dummy[1856], vec_63_bits[57], vec_63_bits[48] );
    foobar f1857( dummy[1857], vec_63_bits[58], vec_63_bits[48] );
    foobar f1858( dummy[1858], vec_63_bits[59], vec_63_bits[48] );
    foobar f1859( dummy[1859], vec_63_bits[60], vec_63_bits[48] );
    foobar f1860( dummy[1860], vec_63_bits[61], vec_63_bits[48] );
    foobar f1861( dummy[1861], vec_63_bits[62], vec_63_bits[48] );
    AN64   an48( o[48], {dummy[1848], dummy[1849], dummy[1850], dummy[1851], dummy[1852], dummy[1853], dummy[1854], dummy[1855], dummy[1856], dummy[1857], dummy[1858], dummy[1859], dummy[1860], dummy[1861], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1862( dummy[1862], vec_63_bits[50], vec_63_bits[49] );
    foobar f1863( dummy[1863], vec_63_bits[51], vec_63_bits[49] );
    foobar f1864( dummy[1864], vec_63_bits[52], vec_63_bits[49] );
    foobar f1865( dummy[1865], vec_63_bits[53], vec_63_bits[49] );
    foobar f1866( dummy[1866], vec_63_bits[54], vec_63_bits[49] );
    foobar f1867( dummy[1867], vec_63_bits[55], vec_63_bits[49] );
    foobar f1868( dummy[1868], vec_63_bits[56], vec_63_bits[49] );
    foobar f1869( dummy[1869], vec_63_bits[57], vec_63_bits[49] );
    foobar f1870( dummy[1870], vec_63_bits[58], vec_63_bits[49] );
    foobar f1871( dummy[1871], vec_63_bits[59], vec_63_bits[49] );
    foobar f1872( dummy[1872], vec_63_bits[60], vec_63_bits[49] );
    foobar f1873( dummy[1873], vec_63_bits[61], vec_63_bits[49] );
    foobar f1874( dummy[1874], vec_63_bits[62], vec_63_bits[49] );
    AN64   an49( o[49], {dummy[1862], dummy[1863], dummy[1864], dummy[1865], dummy[1866], dummy[1867], dummy[1868], dummy[1869], dummy[1870], dummy[1871], dummy[1872], dummy[1873], dummy[1874], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1875( dummy[1875], vec_63_bits[51], vec_63_bits[50] );
    foobar f1876( dummy[1876], vec_63_bits[52], vec_63_bits[50] );
    foobar f1877( dummy[1877], vec_63_bits[53], vec_63_bits[50] );
    foobar f1878( dummy[1878], vec_63_bits[54], vec_63_bits[50] );
    foobar f1879( dummy[1879], vec_63_bits[55], vec_63_bits[50] );
    foobar f1880( dummy[1880], vec_63_bits[56], vec_63_bits[50] );
    foobar f1881( dummy[1881], vec_63_bits[57], vec_63_bits[50] );
    foobar f1882( dummy[1882], vec_63_bits[58], vec_63_bits[50] );
    foobar f1883( dummy[1883], vec_63_bits[59], vec_63_bits[50] );
    foobar f1884( dummy[1884], vec_63_bits[60], vec_63_bits[50] );
    foobar f1885( dummy[1885], vec_63_bits[61], vec_63_bits[50] );
    foobar f1886( dummy[1886], vec_63_bits[62], vec_63_bits[50] );
    AN64   an50( o[50], {dummy[1875], dummy[1876], dummy[1877], dummy[1878], dummy[1879], dummy[1880], dummy[1881], dummy[1882], dummy[1883], dummy[1884], dummy[1885], dummy[1886], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1887( dummy[1887], vec_63_bits[52], vec_63_bits[51] );
    foobar f1888( dummy[1888], vec_63_bits[53], vec_63_bits[51] );
    foobar f1889( dummy[1889], vec_63_bits[54], vec_63_bits[51] );
    foobar f1890( dummy[1890], vec_63_bits[55], vec_63_bits[51] );
    foobar f1891( dummy[1891], vec_63_bits[56], vec_63_bits[51] );
    foobar f1892( dummy[1892], vec_63_bits[57], vec_63_bits[51] );
    foobar f1893( dummy[1893], vec_63_bits[58], vec_63_bits[51] );
    foobar f1894( dummy[1894], vec_63_bits[59], vec_63_bits[51] );
    foobar f1895( dummy[1895], vec_63_bits[60], vec_63_bits[51] );
    foobar f1896( dummy[1896], vec_63_bits[61], vec_63_bits[51] );
    foobar f1897( dummy[1897], vec_63_bits[62], vec_63_bits[51] );
    AN64   an51( o[51], {dummy[1887], dummy[1888], dummy[1889], dummy[1890], dummy[1891], dummy[1892], dummy[1893], dummy[1894], dummy[1895], dummy[1896], dummy[1897], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1898( dummy[1898], vec_63_bits[53], vec_63_bits[52] );
    foobar f1899( dummy[1899], vec_63_bits[54], vec_63_bits[52] );
    foobar f1900( dummy[1900], vec_63_bits[55], vec_63_bits[52] );
    foobar f1901( dummy[1901], vec_63_bits[56], vec_63_bits[52] );
    foobar f1902( dummy[1902], vec_63_bits[57], vec_63_bits[52] );
    foobar f1903( dummy[1903], vec_63_bits[58], vec_63_bits[52] );
    foobar f1904( dummy[1904], vec_63_bits[59], vec_63_bits[52] );
    foobar f1905( dummy[1905], vec_63_bits[60], vec_63_bits[52] );
    foobar f1906( dummy[1906], vec_63_bits[61], vec_63_bits[52] );
    foobar f1907( dummy[1907], vec_63_bits[62], vec_63_bits[52] );
    AN64   an52( o[52], {dummy[1898], dummy[1899], dummy[1900], dummy[1901], dummy[1902], dummy[1903], dummy[1904], dummy[1905], dummy[1906], dummy[1907], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1908( dummy[1908], vec_63_bits[54], vec_63_bits[53] );
    foobar f1909( dummy[1909], vec_63_bits[55], vec_63_bits[53] );
    foobar f1910( dummy[1910], vec_63_bits[56], vec_63_bits[53] );
    foobar f1911( dummy[1911], vec_63_bits[57], vec_63_bits[53] );
    foobar f1912( dummy[1912], vec_63_bits[58], vec_63_bits[53] );
    foobar f1913( dummy[1913], vec_63_bits[59], vec_63_bits[53] );
    foobar f1914( dummy[1914], vec_63_bits[60], vec_63_bits[53] );
    foobar f1915( dummy[1915], vec_63_bits[61], vec_63_bits[53] );
    foobar f1916( dummy[1916], vec_63_bits[62], vec_63_bits[53] );
    AN64   an53( o[53], {dummy[1908], dummy[1909], dummy[1910], dummy[1911], dummy[1912], dummy[1913], dummy[1914], dummy[1915], dummy[1916], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1917( dummy[1917], vec_63_bits[55], vec_63_bits[54] );
    foobar f1918( dummy[1918], vec_63_bits[56], vec_63_bits[54] );
    foobar f1919( dummy[1919], vec_63_bits[57], vec_63_bits[54] );
    foobar f1920( dummy[1920], vec_63_bits[58], vec_63_bits[54] );
    foobar f1921( dummy[1921], vec_63_bits[59], vec_63_bits[54] );
    foobar f1922( dummy[1922], vec_63_bits[60], vec_63_bits[54] );
    foobar f1923( dummy[1923], vec_63_bits[61], vec_63_bits[54] );
    foobar f1924( dummy[1924], vec_63_bits[62], vec_63_bits[54] );
    AN64   an54( o[54], {dummy[1917], dummy[1918], dummy[1919], dummy[1920], dummy[1921], dummy[1922], dummy[1923], dummy[1924], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1925( dummy[1925], vec_63_bits[56], vec_63_bits[55] );
    foobar f1926( dummy[1926], vec_63_bits[57], vec_63_bits[55] );
    foobar f1927( dummy[1927], vec_63_bits[58], vec_63_bits[55] );
    foobar f1928( dummy[1928], vec_63_bits[59], vec_63_bits[55] );
    foobar f1929( dummy[1929], vec_63_bits[60], vec_63_bits[55] );
    foobar f1930( dummy[1930], vec_63_bits[61], vec_63_bits[55] );
    foobar f1931( dummy[1931], vec_63_bits[62], vec_63_bits[55] );
    AN64   an55( o[55], {dummy[1925], dummy[1926], dummy[1927], dummy[1928], dummy[1929], dummy[1930], dummy[1931], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1932( dummy[1932], vec_63_bits[57], vec_63_bits[56] );
    foobar f1933( dummy[1933], vec_63_bits[58], vec_63_bits[56] );
    foobar f1934( dummy[1934], vec_63_bits[59], vec_63_bits[56] );
    foobar f1935( dummy[1935], vec_63_bits[60], vec_63_bits[56] );
    foobar f1936( dummy[1936], vec_63_bits[61], vec_63_bits[56] );
    foobar f1937( dummy[1937], vec_63_bits[62], vec_63_bits[56] );
    AN64   an56( o[56], {dummy[1932], dummy[1933], dummy[1934], dummy[1935], dummy[1936], dummy[1937], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1938( dummy[1938], vec_63_bits[58], vec_63_bits[57] );
    foobar f1939( dummy[1939], vec_63_bits[59], vec_63_bits[57] );
    foobar f1940( dummy[1940], vec_63_bits[60], vec_63_bits[57] );
    foobar f1941( dummy[1941], vec_63_bits[61], vec_63_bits[57] );
    foobar f1942( dummy[1942], vec_63_bits[62], vec_63_bits[57] );
    AN64   an57( o[57], {dummy[1938], dummy[1939], dummy[1940], dummy[1941], dummy[1942], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1943( dummy[1943], vec_63_bits[59], vec_63_bits[58] );
    foobar f1944( dummy[1944], vec_63_bits[60], vec_63_bits[58] );
    foobar f1945( dummy[1945], vec_63_bits[61], vec_63_bits[58] );
    foobar f1946( dummy[1946], vec_63_bits[62], vec_63_bits[58] );
    AN64   an58( o[58], {dummy[1943], dummy[1944], dummy[1945], dummy[1946], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1947( dummy[1947], vec_63_bits[60], vec_63_bits[59] );
    foobar f1948( dummy[1948], vec_63_bits[61], vec_63_bits[59] );
    foobar f1949( dummy[1949], vec_63_bits[62], vec_63_bits[59] );
    AN64   an59( o[59], {dummy[1947], dummy[1948], dummy[1949], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1950( dummy[1950], vec_63_bits[61], vec_63_bits[60] );
    foobar f1951( dummy[1951], vec_63_bits[62], vec_63_bits[60] );
    AN64   an60( o[60], {dummy[1950], dummy[1951], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    foobar f1952( dummy[1952], vec_63_bits[62], vec_63_bits[61] );
    AN64   an61( o[61], {dummy[1952], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
    AN64   an62( o[62], {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } );
endmodule

module gravity_DECoder( o, A, B, C, D, E, F );
    output [62:0] o;
    input A, B, C, D, E, F;
    `wires_2_6
    `wires_3_6
    `wires_4_6
    `wires_5_6
    `wires_6_6
    OR6    o0(  o[0],  A, B, C, D, E, F );
    OR5    o1(  o[1],  E, D, C, B, A );
    OR5    o2(  o[2],  D, C, B, A, EF );
    OR4    o3(  o[3],  D, C, B, A );
    OR5    o4(  o[4],  C, B, A, DF, DE );
    OR4    o5(  o[5],  C, B, A, DE );
    OR4    o6(  o[6],  C, B, A, DEF );
    OR3    o7(  o[7],  C, B, A );
    OR5    o8(  o[8],  B, A, CF, CE, CD );
    OR4    o9(  o[9],  B, A, CE, CD );
    OR4    o10( o[10], B, A, CD, CEF );
    OR3    o11( o[11], B, A, CD );
    OR4    o12( o[12], B, A, CDF, CDE );
    OR3    o13( o[13], B, A, CDE );
    OR3    o14( o[14], B, A, CDEF );
    OR2    o15( o[15], B, A );
    OR5    o16( o[16], A, BF, BE, BD, BC );
    OR4    o17( o[17], A, BE, BD, BC );
    OR4    o18( o[18], A, BD, BC, BEF );
    OR3    o19( o[19], A, BD, BC );
    OR4    o20( o[20], A, BC, BDF, BDE );
    OR3    o21( o[21], A, BC, BDE );
    OR3    o22( o[22], A, BC, BDEF );
    OR2    o23( o[23], A, BC );
    OR4    o24( o[24], A, BCF, BCE, BCD );
    OR3    o25( o[25], A, BCE, BCD );
    OR3    o26( o[26], A, BCD, BCEF );
    OR2    o27( o[27], A, BCD );
    OR3    o28( o[28], A, BCDF, BCDE );
    OR2    o29( o[29], A, BCDE );
    OR2    o30( o[30], A, BCDEF );
    DRIVER o31( o[31], A );
    OR5    o32( o[32], AF, AE, AD, AC, AB );
    OR4    o33( o[33], AE, AD, AC, AB );
    OR4    o34( o[34], AD, AC, AB, AEF );
    OR3    o35( o[35], AD, AC, AB );
    OR4    o36( o[36], AC, AB, ADF, ADE );
    OR3    o37( o[37], AC, AB, ADE );
    OR3    o38( o[38], AC, AB, ADEF );
    OR2    o39( o[39], AC, AB );
    OR4    o40( o[40], AB, ACF, ACE, ACD );
    OR3    o41( o[41], AB, ACE, ACD );
    OR3    o42( o[42], AB, ACD, ACEF );
    OR2    o43( o[43], AB, ACD );
    OR3    o44( o[44], AB, ACDF, ACDE );
    OR2    o45( o[45], AB, ACDE );
    OR2    o46( o[46], AB, ACDEF );
    DRIVER o47( o[47], AB );
    OR4    o48( o[48], ABF, ABE, ABD, ABC );
    OR3    o49( o[49], ABE, ABD, ABC );
    OR3    o50( o[50], ABD, ABC, ABEF );
    OR2    o51( o[51], ABD, ABC );
    OR3    o52( o[52], ABC, ABDF, ABDE );
    OR2    o53( o[53], ABC, ABDE );
    OR2    o54( o[54], ABC, ABDEF );
    DRIVER o55( o[55], ABC );
    OR3    o56( o[56], ABCF, ABCE, ABCD );
    OR2    o57( o[57], ABCE, ABCD );
    OR2    o58( o[58], ABCD, ABCEF );
    DRIVER o59( o[59], ABCD );
    OR2    o60( o[60], ABCDF, ABCDE );
    DRIVER o61( o[61], ABCDE );
    DRIVER o62( o[62], ABCDEF );
endmodule

module THRES_1_5( o, A, B, C, D, E );
    input  A, B, C, D, E;
    output o;
    OR5  ret( o, A, B, C, D, E );
endmodule

module THRES_2_5( o, A, B, C, D, E );
    input  A, B, C, D, E;
    output o;
    `wires_2_5
    OR15 ret( o, {AB, AC, AD, AE, BC, BD, BE, CD, CE, DE} );
endmodule

module THRES_3_5( o, A, B, C, D, E );
    input  A, B, C, D, E;
    output o;
    `wires_3_5
    OR20 ret( o, {ABC, ABD, ABE, ACD, ACE, ADE, BCD, BCE, BDE, CDE} );
endmodule

module THRES_4_5( o, A, B, C, D, E );
    input  A, B, C, D, E;
    output o;
    `wires_4_5
    OR15 ret( o, {ABCD, ABCE, ABDE, ACDE, BCDE} );
endmodule

module THRES_5_5( o, A, B, C, D, E );
    input  A, B, C, D, E;
    output o;
    `wires_5_5
    DRIVER ret( o, ABCDE );
endmodule

module gravity_ENCoder( o, i );
    inout      [62:0]   i;
    output     [ 5:0]   o;
    wire       [62:0]   I;

    Sanitizer s(I, i);

    OR32 o0( o[0], {
        I[0],  I[2],  I[4],  I[6],  I[8],  I[10], I[12], I[14],
        I[16], I[18], I[20], I[22], I[24], I[26], I[28], I[30],
        I[32], I[34], I[36], I[38], I[40], I[42], I[44], I[46],
        I[48], I[50], I[52], I[54], I[56], I[58], I[60], I[62]
        } );
    OR32 o1( o[1], {
       I[1],  I[2],  I[5],  I[6],  I[9],  I[10], I[13], I[14],
       I[17], I[18], I[21], I[22], I[25], I[26], I[29], I[30],
       I[33], I[34], I[37], I[38], I[41], I[42], I[45], I[46],
       I[49], I[50], I[53], I[54], I[57], I[58], I[61], I[62]
       } );
    OR32 o2( o[2], {
       I[3],  I[4],  I[5],  I[6],  I[11], I[12], I[13], I[14],
       I[19], I[20], I[21], I[22], I[27], I[28], I[29], I[30],
       I[35], I[36], I[37], I[38], I[43], I[44], I[45], I[46],
       I[51], I[52], I[53], I[54], I[59], I[60], I[61], I[62]
       } );
    OR32 o3( o[3], {
       I[7],  I[8],  I[9],  I[10], I[11], I[12], I[13], I[14],
       I[23], I[24], I[25], I[26], I[27], I[28], I[29], I[30],
       I[39], I[40], I[41], I[42], I[43], I[44], I[45], I[46],
       I[55], I[56], I[57], I[58], I[59], I[60], I[61], I[62]
       } );
    OR32 o4( o[4], {
       I[15], I[16], I[17], I[18], I[19], I[20], I[21], I[22],
       I[23], I[24], I[25], I[26], I[27], I[28], I[29], I[30],
       I[47], I[48], I[49], I[50], I[51], I[52], I[53], I[54],
       I[55], I[56], I[57], I[58], I[59], I[60], I[61], I[62]
       } );
    OR32 o5( o[5], {
       I[31], I[32], I[33], I[34], I[35], I[36], I[37], I[38],
       I[39], I[40], I[41], I[42], I[43], I[44], I[45], I[46],
       I[47], I[48], I[49], I[50], I[51], I[52], I[53], I[54],
       I[55], I[56], I[57], I[58], I[59], I[60], I[61], I[62]
       } );

endmodule

module THRES_1_5_VEC( o, A, B, C, D, E );
    THRES_1_5 t00( o[0],  A[0],  B[0],  C[0],  D[0],  E[0] );
    THRES_1_5 t01( o[1],  A[1],  B[1],  C[1],  D[1],  E[1] );
    THRES_1_5 t02( o[2],  A[2],  B[2],  C[2],  D[2],  E[2] );
    THRES_1_5 t03( o[3],  A[3],  B[3],  C[3],  D[3],  E[3] );
    THRES_1_5 t04( o[4],  A[4],  B[4],  C[4],  D[4],  E[4] );
    THRES_1_5 t05( o[5],  A[5],  B[5],  C[5],  D[5],  E[5] );
    THRES_1_5 t06( o[6],  A[6],  B[6],  C[6],  D[6],  E[6] );
    THRES_1_5 t07( o[7],  A[7],  B[7],  C[7],  D[7],  E[7] );
    THRES_1_5 t08( o[8],  A[8],  B[8],  C[8],  D[8],  E[8] );
    THRES_1_5 t09( o[9],  A[9],  B[9],  C[9],  D[9],  E[9] );
    THRES_1_5 t10( o[10], A[10], B[10], C[10], D[10], E[10] );
    THRES_1_5 t11( o[11], A[11], B[11], C[11], D[11], E[11] );
    THRES_1_5 t12( o[12], A[12], B[12], C[12], D[12], E[12] );
    THRES_1_5 t13( o[13], A[13], B[13], C[13], D[13], E[13] );
    THRES_1_5 t14( o[14], A[14], B[14], C[14], D[14], E[14] );
    THRES_1_5 t15( o[15], A[15], B[15], C[15], D[15], E[15] );
    THRES_1_5 t16( o[16], A[16], B[16], C[16], D[16], E[16] );
    THRES_1_5 t17( o[17], A[17], B[17], C[17], D[17], E[17] );
    THRES_1_5 t18( o[18], A[18], B[18], C[18], D[18], E[18] );
    THRES_1_5 t19( o[19], A[19], B[19], C[19], D[19], E[19] );
    THRES_1_5 t20( o[20], A[20], B[20], C[20], D[20], E[20] );
    THRES_1_5 t21( o[21], A[21], B[21], C[21], D[21], E[21] );
    THRES_1_5 t22( o[22], A[22], B[22], C[22], D[22], E[22] );
    THRES_1_5 t23( o[23], A[23], B[23], C[23], D[23], E[23] );
    THRES_1_5 t24( o[24], A[24], B[24], C[24], D[24], E[24] );
    THRES_1_5 t25( o[25], A[25], B[25], C[25], D[25], E[25] );
    THRES_1_5 t26( o[26], A[26], B[26], C[26], D[26], E[26] );
    THRES_1_5 t27( o[27], A[27], B[27], C[27], D[27], E[27] );
    THRES_1_5 t28( o[28], A[28], B[28], C[28], D[28], E[28] );
    THRES_1_5 t29( o[29], A[29], B[29], C[29], D[29], E[29] );
    THRES_1_5 t30( o[30], A[30], B[30], C[30], D[30], E[30] );
    THRES_1_5 t31( o[31], A[31], B[31], C[31], D[31], E[31] );
    THRES_1_5 t32( o[32], A[32], B[32], C[32], D[32], E[32] );
    THRES_1_5 t33( o[33], A[33], B[33], C[33], D[33], E[33] );
    THRES_1_5 t34( o[34], A[34], B[34], C[34], D[34], E[34] );
    THRES_1_5 t35( o[35], A[35], B[35], C[35], D[35], E[35] );
    THRES_1_5 t36( o[36], A[36], B[36], C[36], D[36], E[36] );
    THRES_1_5 t37( o[37], A[37], B[37], C[37], D[37], E[37] );
    THRES_1_5 t38( o[38], A[38], B[38], C[38], D[38], E[38] );
    THRES_1_5 t39( o[39], A[39], B[39], C[39], D[39], E[39] );
    THRES_1_5 t40( o[40], A[40], B[40], C[40], D[40], E[40] );
    THRES_1_5 t41( o[41], A[41], B[41], C[41], D[41], E[41] );
    THRES_1_5 t42( o[42], A[42], B[42], C[42], D[42], E[42] );
    THRES_1_5 t43( o[43], A[43], B[43], C[43], D[43], E[43] );
    THRES_1_5 t44( o[44], A[44], B[44], C[44], D[44], E[44] );
    THRES_1_5 t45( o[45], A[45], B[45], C[45], D[45], E[45] );
    THRES_1_5 t46( o[46], A[46], B[46], C[46], D[46], E[46] );
    THRES_1_5 t47( o[47], A[47], B[47], C[47], D[47], E[47] );
    THRES_1_5 t48( o[48], A[48], B[48], C[48], D[48], E[48] );
    THRES_1_5 t49( o[49], A[49], B[49], C[49], D[49], E[49] );
    THRES_1_5 t50( o[50], A[50], B[50], C[50], D[50], E[50] );
    THRES_1_5 t51( o[51], A[51], B[51], C[51], D[51], E[51] );
    THRES_1_5 t52( o[52], A[52], B[52], C[52], D[52], E[52] );
    THRES_1_5 t53( o[53], A[53], B[53], C[53], D[53], E[53] );
    THRES_1_5 t54( o[54], A[54], B[54], C[54], D[54], E[54] );
    THRES_1_5 t55( o[55], A[55], B[55], C[55], D[55], E[55] );
    THRES_1_5 t56( o[56], A[56], B[56], C[56], D[56], E[56] );
    THRES_1_5 t57( o[57], A[57], B[57], C[57], D[57], E[57] );
    THRES_1_5 t58( o[58], A[58], B[58], C[58], D[58], E[58] );
    THRES_1_5 t59( o[59], A[59], B[59], C[59], D[59], E[59] );
    THRES_1_5 t60( o[60], A[60], B[60], C[60], D[60], E[60] );
    THRES_1_5 t61( o[61], A[61], B[61], C[61], D[61], E[61] );
    THRES_1_5 t62( o[62], A[62], B[62], C[62], D[62], E[62] );
endmodule

module THRES_2_5_VEC( o, A, B, C, D, E );
    THRES_2_5 t00( o[0],  A[0],  B[0],  C[0],  D[0],  E[0] );
    THRES_2_5 t01( o[1],  A[1],  B[1],  C[1],  D[1],  E[1] );
    THRES_2_5 t02( o[2],  A[2],  B[2],  C[2],  D[2],  E[2] );
    THRES_2_5 t03( o[3],  A[3],  B[3],  C[3],  D[3],  E[3] );
    THRES_2_5 t04( o[4],  A[4],  B[4],  C[4],  D[4],  E[4] );
    THRES_2_5 t05( o[5],  A[5],  B[5],  C[5],  D[5],  E[5] );
    THRES_2_5 t06( o[6],  A[6],  B[6],  C[6],  D[6],  E[6] );
    THRES_2_5 t07( o[7],  A[7],  B[7],  C[7],  D[7],  E[7] );
    THRES_2_5 t08( o[8],  A[8],  B[8],  C[8],  D[8],  E[8] );
    THRES_2_5 t09( o[9],  A[9],  B[9],  C[9],  D[9],  E[9] );
    THRES_2_5 t10( o[10], A[10], B[10], C[10], D[10], E[10] );
    THRES_2_5 t11( o[11], A[11], B[11], C[11], D[11], E[11] );
    THRES_2_5 t12( o[12], A[12], B[12], C[12], D[12], E[12] );
    THRES_2_5 t13( o[13], A[13], B[13], C[13], D[13], E[13] );
    THRES_2_5 t14( o[14], A[14], B[14], C[14], D[14], E[14] );
    THRES_2_5 t15( o[15], A[15], B[15], C[15], D[15], E[15] );
    THRES_2_5 t16( o[16], A[16], B[16], C[16], D[16], E[16] );
    THRES_2_5 t17( o[17], A[17], B[17], C[17], D[17], E[17] );
    THRES_2_5 t18( o[18], A[18], B[18], C[18], D[18], E[18] );
    THRES_2_5 t19( o[19], A[19], B[19], C[19], D[19], E[19] );
    THRES_2_5 t20( o[20], A[20], B[20], C[20], D[20], E[20] );
    THRES_2_5 t21( o[21], A[21], B[21], C[21], D[21], E[21] );
    THRES_2_5 t22( o[22], A[22], B[22], C[22], D[22], E[22] );
    THRES_2_5 t23( o[23], A[23], B[23], C[23], D[23], E[23] );
    THRES_2_5 t24( o[24], A[24], B[24], C[24], D[24], E[24] );
    THRES_2_5 t25( o[25], A[25], B[25], C[25], D[25], E[25] );
    THRES_2_5 t26( o[26], A[26], B[26], C[26], D[26], E[26] );
    THRES_2_5 t27( o[27], A[27], B[27], C[27], D[27], E[27] );
    THRES_2_5 t28( o[28], A[28], B[28], C[28], D[28], E[28] );
    THRES_2_5 t29( o[29], A[29], B[29], C[29], D[29], E[29] );
    THRES_2_5 t30( o[30], A[30], B[30], C[30], D[30], E[30] );
    THRES_2_5 t31( o[31], A[31], B[31], C[31], D[31], E[31] );
    THRES_2_5 t32( o[32], A[32], B[32], C[32], D[32], E[32] );
    THRES_2_5 t33( o[33], A[33], B[33], C[33], D[33], E[33] );
    THRES_2_5 t34( o[34], A[34], B[34], C[34], D[34], E[34] );
    THRES_2_5 t35( o[35], A[35], B[35], C[35], D[35], E[35] );
    THRES_2_5 t36( o[36], A[36], B[36], C[36], D[36], E[36] );
    THRES_2_5 t37( o[37], A[37], B[37], C[37], D[37], E[37] );
    THRES_2_5 t38( o[38], A[38], B[38], C[38], D[38], E[38] );
    THRES_2_5 t39( o[39], A[39], B[39], C[39], D[39], E[39] );
    THRES_2_5 t40( o[40], A[40], B[40], C[40], D[40], E[40] );
    THRES_2_5 t41( o[41], A[41], B[41], C[41], D[41], E[41] );
    THRES_2_5 t42( o[42], A[42], B[42], C[42], D[42], E[42] );
    THRES_2_5 t43( o[43], A[43], B[43], C[43], D[43], E[43] );
    THRES_2_5 t44( o[44], A[44], B[44], C[44], D[44], E[44] );
    THRES_2_5 t45( o[45], A[45], B[45], C[45], D[45], E[45] );
    THRES_2_5 t46( o[46], A[46], B[46], C[46], D[46], E[46] );
    THRES_2_5 t47( o[47], A[47], B[47], C[47], D[47], E[47] );
    THRES_2_5 t48( o[48], A[48], B[48], C[48], D[48], E[48] );
    THRES_2_5 t49( o[49], A[49], B[49], C[49], D[49], E[49] );
    THRES_2_5 t50( o[50], A[50], B[50], C[50], D[50], E[50] );
    THRES_2_5 t51( o[51], A[51], B[51], C[51], D[51], E[51] );
    THRES_2_5 t52( o[52], A[52], B[52], C[52], D[52], E[52] );
    THRES_2_5 t53( o[53], A[53], B[53], C[53], D[53], E[53] );
    THRES_2_5 t54( o[54], A[54], B[54], C[54], D[54], E[54] );
    THRES_2_5 t55( o[55], A[55], B[55], C[55], D[55], E[55] );
    THRES_2_5 t56( o[56], A[56], B[56], C[56], D[56], E[56] );
    THRES_2_5 t57( o[57], A[57], B[57], C[57], D[57], E[57] );
    THRES_2_5 t58( o[58], A[58], B[58], C[58], D[58], E[58] );
    THRES_2_5 t59( o[59], A[59], B[59], C[59], D[59], E[59] );
    THRES_2_5 t60( o[60], A[60], B[60], C[60], D[60], E[60] );
    THRES_2_5 t61( o[61], A[61], B[61], C[61], D[61], E[61] );
    THRES_2_5 t62( o[62], A[62], B[62], C[62], D[62], E[62] );
endmodule

module THRES_3_5_VEC( o, A, B, C, D, E );
    THRES_3_5 t00( o[0],  A[0],  B[0],  C[0],  D[0],  E[0] );
    THRES_3_5 t01( o[1],  A[1],  B[1],  C[1],  D[1],  E[1] );
    THRES_3_5 t02( o[2],  A[2],  B[2],  C[2],  D[2],  E[2] );
    THRES_3_5 t03( o[3],  A[3],  B[3],  C[3],  D[3],  E[3] );
    THRES_3_5 t04( o[4],  A[4],  B[4],  C[4],  D[4],  E[4] );
    THRES_3_5 t05( o[5],  A[5],  B[5],  C[5],  D[5],  E[5] );
    THRES_3_5 t06( o[6],  A[6],  B[6],  C[6],  D[6],  E[6] );
    THRES_3_5 t07( o[7],  A[7],  B[7],  C[7],  D[7],  E[7] );
    THRES_3_5 t08( o[8],  A[8],  B[8],  C[8],  D[8],  E[8] );
    THRES_3_5 t09( o[9],  A[9],  B[9],  C[9],  D[9],  E[9] );
    THRES_3_5 t10( o[10], A[10], B[10], C[10], D[10], E[10] );
    THRES_3_5 t11( o[11], A[11], B[11], C[11], D[11], E[11] );
    THRES_3_5 t12( o[12], A[12], B[12], C[12], D[12], E[12] );
    THRES_3_5 t13( o[13], A[13], B[13], C[13], D[13], E[13] );
    THRES_3_5 t14( o[14], A[14], B[14], C[14], D[14], E[14] );
    THRES_3_5 t15( o[15], A[15], B[15], C[15], D[15], E[15] );
    THRES_3_5 t16( o[16], A[16], B[16], C[16], D[16], E[16] );
    THRES_3_5 t17( o[17], A[17], B[17], C[17], D[17], E[17] );
    THRES_3_5 t18( o[18], A[18], B[18], C[18], D[18], E[18] );
    THRES_3_5 t19( o[19], A[19], B[19], C[19], D[19], E[19] );
    THRES_3_5 t20( o[20], A[20], B[20], C[20], D[20], E[20] );
    THRES_3_5 t21( o[21], A[21], B[21], C[21], D[21], E[21] );
    THRES_3_5 t22( o[22], A[22], B[22], C[22], D[22], E[22] );
    THRES_3_5 t23( o[23], A[23], B[23], C[23], D[23], E[23] );
    THRES_3_5 t24( o[24], A[24], B[24], C[24], D[24], E[24] );
    THRES_3_5 t25( o[25], A[25], B[25], C[25], D[25], E[25] );
    THRES_3_5 t26( o[26], A[26], B[26], C[26], D[26], E[26] );
    THRES_3_5 t27( o[27], A[27], B[27], C[27], D[27], E[27] );
    THRES_3_5 t28( o[28], A[28], B[28], C[28], D[28], E[28] );
    THRES_3_5 t29( o[29], A[29], B[29], C[29], D[29], E[29] );
    THRES_3_5 t30( o[30], A[30], B[30], C[30], D[30], E[30] );
    THRES_3_5 t31( o[31], A[31], B[31], C[31], D[31], E[31] );
    THRES_3_5 t32( o[32], A[32], B[32], C[32], D[32], E[32] );
    THRES_3_5 t33( o[33], A[33], B[33], C[33], D[33], E[33] );
    THRES_3_5 t34( o[34], A[34], B[34], C[34], D[34], E[34] );
    THRES_3_5 t35( o[35], A[35], B[35], C[35], D[35], E[35] );
    THRES_3_5 t36( o[36], A[36], B[36], C[36], D[36], E[36] );
    THRES_3_5 t37( o[37], A[37], B[37], C[37], D[37], E[37] );
    THRES_3_5 t38( o[38], A[38], B[38], C[38], D[38], E[38] );
    THRES_3_5 t39( o[39], A[39], B[39], C[39], D[39], E[39] );
    THRES_3_5 t40( o[40], A[40], B[40], C[40], D[40], E[40] );
    THRES_3_5 t41( o[41], A[41], B[41], C[41], D[41], E[41] );
    THRES_3_5 t42( o[42], A[42], B[42], C[42], D[42], E[42] );
    THRES_3_5 t43( o[43], A[43], B[43], C[43], D[43], E[43] );
    THRES_3_5 t44( o[44], A[44], B[44], C[44], D[44], E[44] );
    THRES_3_5 t45( o[45], A[45], B[45], C[45], D[45], E[45] );
    THRES_3_5 t46( o[46], A[46], B[46], C[46], D[46], E[46] );
    THRES_3_5 t47( o[47], A[47], B[47], C[47], D[47], E[47] );
    THRES_3_5 t48( o[48], A[48], B[48], C[48], D[48], E[48] );
    THRES_3_5 t49( o[49], A[49], B[49], C[49], D[49], E[49] );
    THRES_3_5 t50( o[50], A[50], B[50], C[50], D[50], E[50] );
    THRES_3_5 t51( o[51], A[51], B[51], C[51], D[51], E[51] );
    THRES_3_5 t52( o[52], A[52], B[52], C[52], D[52], E[52] );
    THRES_3_5 t53( o[53], A[53], B[53], C[53], D[53], E[53] );
    THRES_3_5 t54( o[54], A[54], B[54], C[54], D[54], E[54] );
    THRES_3_5 t55( o[55], A[55], B[55], C[55], D[55], E[55] );
    THRES_3_5 t56( o[56], A[56], B[56], C[56], D[56], E[56] );
    THRES_3_5 t57( o[57], A[57], B[57], C[57], D[57], E[57] );
    THRES_3_5 t58( o[58], A[58], B[58], C[58], D[58], E[58] );
    THRES_3_5 t59( o[59], A[59], B[59], C[59], D[59], E[59] );
    THRES_3_5 t60( o[60], A[60], B[60], C[60], D[60], E[60] );
    THRES_3_5 t61( o[61], A[61], B[61], C[61], D[61], E[61] );
    THRES_3_5 t62( o[62], A[62], B[62], C[62], D[62], E[62] );
endmodule

module THRES_4_5_VEC( o, A, B, C, D, E );
    THRES_4_5 t00( o[0],  A[0],  B[0],  C[0],  D[0],  E[0] );
    THRES_4_5 t01( o[1],  A[1],  B[1],  C[1],  D[1],  E[1] );
    THRES_4_5 t02( o[2],  A[2],  B[2],  C[2],  D[2],  E[2] );
    THRES_4_5 t03( o[3],  A[3],  B[3],  C[3],  D[3],  E[3] );
    THRES_4_5 t04( o[4],  A[4],  B[4],  C[4],  D[4],  E[4] );
    THRES_4_5 t05( o[5],  A[5],  B[5],  C[5],  D[5],  E[5] );
    THRES_4_5 t06( o[6],  A[6],  B[6],  C[6],  D[6],  E[6] );
    THRES_4_5 t07( o[7],  A[7],  B[7],  C[7],  D[7],  E[7] );
    THRES_4_5 t08( o[8],  A[8],  B[8],  C[8],  D[8],  E[8] );
    THRES_4_5 t09( o[9],  A[9],  B[9],  C[9],  D[9],  E[9] );
    THRES_4_5 t10( o[10], A[10], B[10], C[10], D[10], E[10] );
    THRES_4_5 t11( o[11], A[11], B[11], C[11], D[11], E[11] );
    THRES_4_5 t12( o[12], A[12], B[12], C[12], D[12], E[12] );
    THRES_4_5 t13( o[13], A[13], B[13], C[13], D[13], E[13] );
    THRES_4_5 t14( o[14], A[14], B[14], C[14], D[14], E[14] );
    THRES_4_5 t15( o[15], A[15], B[15], C[15], D[15], E[15] );
    THRES_4_5 t16( o[16], A[16], B[16], C[16], D[16], E[16] );
    THRES_4_5 t17( o[17], A[17], B[17], C[17], D[17], E[17] );
    THRES_4_5 t18( o[18], A[18], B[18], C[18], D[18], E[18] );
    THRES_4_5 t19( o[19], A[19], B[19], C[19], D[19], E[19] );
    THRES_4_5 t20( o[20], A[20], B[20], C[20], D[20], E[20] );
    THRES_4_5 t21( o[21], A[21], B[21], C[21], D[21], E[21] );
    THRES_4_5 t22( o[22], A[22], B[22], C[22], D[22], E[22] );
    THRES_4_5 t23( o[23], A[23], B[23], C[23], D[23], E[23] );
    THRES_4_5 t24( o[24], A[24], B[24], C[24], D[24], E[24] );
    THRES_4_5 t25( o[25], A[25], B[25], C[25], D[25], E[25] );
    THRES_4_5 t26( o[26], A[26], B[26], C[26], D[26], E[26] );
    THRES_4_5 t27( o[27], A[27], B[27], C[27], D[27], E[27] );
    THRES_4_5 t28( o[28], A[28], B[28], C[28], D[28], E[28] );
    THRES_4_5 t29( o[29], A[29], B[29], C[29], D[29], E[29] );
    THRES_4_5 t30( o[30], A[30], B[30], C[30], D[30], E[30] );
    THRES_4_5 t31( o[31], A[31], B[31], C[31], D[31], E[31] );
    THRES_4_5 t32( o[32], A[32], B[32], C[32], D[32], E[32] );
    THRES_4_5 t33( o[33], A[33], B[33], C[33], D[33], E[33] );
    THRES_4_5 t34( o[34], A[34], B[34], C[34], D[34], E[34] );
    THRES_4_5 t35( o[35], A[35], B[35], C[35], D[35], E[35] );
    THRES_4_5 t36( o[36], A[36], B[36], C[36], D[36], E[36] );
    THRES_4_5 t37( o[37], A[37], B[37], C[37], D[37], E[37] );
    THRES_4_5 t38( o[38], A[38], B[38], C[38], D[38], E[38] );
    THRES_4_5 t39( o[39], A[39], B[39], C[39], D[39], E[39] );
    THRES_4_5 t40( o[40], A[40], B[40], C[40], D[40], E[40] );
    THRES_4_5 t41( o[41], A[41], B[41], C[41], D[41], E[41] );
    THRES_4_5 t42( o[42], A[42], B[42], C[42], D[42], E[42] );
    THRES_4_5 t43( o[43], A[43], B[43], C[43], D[43], E[43] );
    THRES_4_5 t44( o[44], A[44], B[44], C[44], D[44], E[44] );
    THRES_4_5 t45( o[45], A[45], B[45], C[45], D[45], E[45] );
    THRES_4_5 t46( o[46], A[46], B[46], C[46], D[46], E[46] );
    THRES_4_5 t47( o[47], A[47], B[47], C[47], D[47], E[47] );
    THRES_4_5 t48( o[48], A[48], B[48], C[48], D[48], E[48] );
    THRES_4_5 t49( o[49], A[49], B[49], C[49], D[49], E[49] );
    THRES_4_5 t50( o[50], A[50], B[50], C[50], D[50], E[50] );
    THRES_4_5 t51( o[51], A[51], B[51], C[51], D[51], E[51] );
    THRES_4_5 t52( o[52], A[52], B[52], C[52], D[52], E[52] );
    THRES_4_5 t53( o[53], A[53], B[53], C[53], D[53], E[53] );
    THRES_4_5 t54( o[54], A[54], B[54], C[54], D[54], E[54] );
    THRES_4_5 t55( o[55], A[55], B[55], C[55], D[55], E[55] );
    THRES_4_5 t56( o[56], A[56], B[56], C[56], D[56], E[56] );
    THRES_4_5 t57( o[57], A[57], B[57], C[57], D[57], E[57] );
    THRES_4_5 t58( o[58], A[58], B[58], C[58], D[58], E[58] );
    THRES_4_5 t59( o[59], A[59], B[59], C[59], D[59], E[59] );
    THRES_4_5 t60( o[60], A[60], B[60], C[60], D[60], E[60] );
    THRES_4_5 t61( o[61], A[61], B[61], C[61], D[61], E[61] );
    THRES_4_5 t62( o[62], A[62], B[62], C[62], D[62], E[62] );
endmodule

module THRES_5_5_VEC( o, A, B, C, D, E );
    THRES_5_5 t00( o[0],  A[0],  B[0],  C[0],  D[0],  E[0] );
    THRES_5_5 t01( o[1],  A[1],  B[1],  C[1],  D[1],  E[1] );
    THRES_5_5 t02( o[2],  A[2],  B[2],  C[2],  D[2],  E[2] );
    THRES_5_5 t03( o[3],  A[3],  B[3],  C[3],  D[3],  E[3] );
    THRES_5_5 t04( o[4],  A[4],  B[4],  C[4],  D[4],  E[4] );
    THRES_5_5 t05( o[5],  A[5],  B[5],  C[5],  D[5],  E[5] );
    THRES_5_5 t06( o[6],  A[6],  B[6],  C[6],  D[6],  E[6] );
    THRES_5_5 t07( o[7],  A[7],  B[7],  C[7],  D[7],  E[7] );
    THRES_5_5 t08( o[8],  A[8],  B[8],  C[8],  D[8],  E[8] );
    THRES_5_5 t09( o[9],  A[9],  B[9],  C[9],  D[9],  E[9] );
    THRES_5_5 t10( o[10], A[10], B[10], C[10], D[10], E[10] );
    THRES_5_5 t11( o[11], A[11], B[11], C[11], D[11], E[11] );
    THRES_5_5 t12( o[12], A[12], B[12], C[12], D[12], E[12] );
    THRES_5_5 t13( o[13], A[13], B[13], C[13], D[13], E[13] );
    THRES_5_5 t14( o[14], A[14], B[14], C[14], D[14], E[14] );
    THRES_5_5 t15( o[15], A[15], B[15], C[15], D[15], E[15] );
    THRES_5_5 t16( o[16], A[16], B[16], C[16], D[16], E[16] );
    THRES_5_5 t17( o[17], A[17], B[17], C[17], D[17], E[17] );
    THRES_5_5 t18( o[18], A[18], B[18], C[18], D[18], E[18] );
    THRES_5_5 t19( o[19], A[19], B[19], C[19], D[19], E[19] );
    THRES_5_5 t20( o[20], A[20], B[20], C[20], D[20], E[20] );
    THRES_5_5 t21( o[21], A[21], B[21], C[21], D[21], E[21] );
    THRES_5_5 t22( o[22], A[22], B[22], C[22], D[22], E[22] );
    THRES_5_5 t23( o[23], A[23], B[23], C[23], D[23], E[23] );
    THRES_5_5 t24( o[24], A[24], B[24], C[24], D[24], E[24] );
    THRES_5_5 t25( o[25], A[25], B[25], C[25], D[25], E[25] );
    THRES_5_5 t26( o[26], A[26], B[26], C[26], D[26], E[26] );
    THRES_5_5 t27( o[27], A[27], B[27], C[27], D[27], E[27] );
    THRES_5_5 t28( o[28], A[28], B[28], C[28], D[28], E[28] );
    THRES_5_5 t29( o[29], A[29], B[29], C[29], D[29], E[29] );
    THRES_5_5 t30( o[30], A[30], B[30], C[30], D[30], E[30] );
    THRES_5_5 t31( o[31], A[31], B[31], C[31], D[31], E[31] );
    THRES_5_5 t32( o[32], A[32], B[32], C[32], D[32], E[32] );
    THRES_5_5 t33( o[33], A[33], B[33], C[33], D[33], E[33] );
    THRES_5_5 t34( o[34], A[34], B[34], C[34], D[34], E[34] );
    THRES_5_5 t35( o[35], A[35], B[35], C[35], D[35], E[35] );
    THRES_5_5 t36( o[36], A[36], B[36], C[36], D[36], E[36] );
    THRES_5_5 t37( o[37], A[37], B[37], C[37], D[37], E[37] );
    THRES_5_5 t38( o[38], A[38], B[38], C[38], D[38], E[38] );
    THRES_5_5 t39( o[39], A[39], B[39], C[39], D[39], E[39] );
    THRES_5_5 t40( o[40], A[40], B[40], C[40], D[40], E[40] );
    THRES_5_5 t41( o[41], A[41], B[41], C[41], D[41], E[41] );
    THRES_5_5 t42( o[42], A[42], B[42], C[42], D[42], E[42] );
    THRES_5_5 t43( o[43], A[43], B[43], C[43], D[43], E[43] );
    THRES_5_5 t44( o[44], A[44], B[44], C[44], D[44], E[44] );
    THRES_5_5 t45( o[45], A[45], B[45], C[45], D[45], E[45] );
    THRES_5_5 t46( o[46], A[46], B[46], C[46], D[46], E[46] );
    THRES_5_5 t47( o[47], A[47], B[47], C[47], D[47], E[47] );
    THRES_5_5 t48( o[48], A[48], B[48], C[48], D[48], E[48] );
    THRES_5_5 t49( o[49], A[49], B[49], C[49], D[49], E[49] );
    THRES_5_5 t50( o[50], A[50], B[50], C[50], D[50], E[50] );
    THRES_5_5 t51( o[51], A[51], B[51], C[51], D[51], E[51] );
    THRES_5_5 t52( o[52], A[52], B[52], C[52], D[52], E[52] );
    THRES_5_5 t53( o[53], A[53], B[53], C[53], D[53], E[53] );
    THRES_5_5 t54( o[54], A[54], B[54], C[54], D[54], E[54] );
    THRES_5_5 t55( o[55], A[55], B[55], C[55], D[55], E[55] );
    THRES_5_5 t56( o[56], A[56], B[56], C[56], D[56], E[56] );
    THRES_5_5 t57( o[57], A[57], B[57], C[57], D[57], E[57] );
    THRES_5_5 t58( o[58], A[58], B[58], C[58], D[58], E[58] );
    THRES_5_5 t59( o[59], A[59], B[59], C[59], D[59], E[59] );
    THRES_5_5 t60( o[60], A[60], B[60], C[60], D[60], E[60] );
    THRES_5_5 t61( o[61], A[61], B[61], C[61], D[61], E[61] );
    THRES_5_5 t62( o[62], A[62], B[62], C[62], D[62], E[62] );
endmodule

module gravity_SORT(rank0, rank1, rank2, rank3, rank4, i0, i1, i2, i3, i4);
	input  [5:0] i0, i1, i2, i3, i4;
	output [5:0] rank0, rank1, rank2, rank3, rank4;
    wire   [62:0] I0, I1, I2, I3, I4;
    wire   [62:0] w0, w1, w2, w3, w4;
    wire   [62:0] rank0_raw, rank1_raw, rank2_raw, rank3_raw, rank4_raw;

    gravity_DECoder dec_0( I0, i0[5], i0[4], i0[3], i0[2], i0[1], i0[0] );
    gravity_DECoder dec_1( I1, i1[5], i1[4], i1[3], i1[2], i1[1], i1[0] );
    gravity_DECoder dec_2( I2, i2[5], i2[4], i2[3], i2[2], i2[1], i2[0] );
    gravity_DECoder dec_3( I3, i3[5], i3[4], i3[3], i3[2], i3[1], i3[0] );
    gravity_DECoder dec_4( I4, i4[5], i4[4], i4[3], i4[2], i4[1], i4[0] );

    THRES_1_5       thres_rank0_raw [62:0]( w0, I0, I1, I2, I3, I4);
    THRES_2_5       thres_rank1_raw [62:0]( w1, I0, I1, I2, I3, I4);
    THRES_3_5       thres_rank2_raw [62:0]( w2, I0, I1, I2, I3, I4);
    THRES_4_5       thres_rank3_raw [62:0]( w3, I0, I1, I2, I3, I4);
    THRES_5_5       thres_rank4_raw [62:0]( w4, I0, I1, I2, I3, I4);

    gravity_ENCoder result0( rank0, w0 );
    gravity_ENCoder result1( rank1, w1 );
    gravity_ENCoder result2( rank2, w2 );
    gravity_ENCoder result3( rank3, w3 );
    gravity_ENCoder result4( rank4, w4 );

endmodule

module sorting(rank0, rank1, rank2, rank3, rank4, i0, i1, i2, i3, i4);
//DO NOT CHANGE!
	input  [5:0] i0, i1, i2, i3, i4;
	output [5:0] rank0, rank1, rank2, rank3, rank4;
//---------------------------------------------------
    gravity_SORT Newton(
        rank0, rank1, rank2, rank3, rank4,
        i0, i1, i2, i3, i4
    );

endmodule
